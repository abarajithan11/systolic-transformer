##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Thu Mar 23 02:03:03 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO dualcore
  CLASS BLOCK ;
  SIZE 546.600000 BY 545.600000 ;
  FOREIGN dualcore 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 231.300000 0.600000 231.500000 ;
    END
  END clk1
  PIN rst1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 234.500000 0.600000 234.700000 ;
    END
  END rst1
  PIN mem_in_core1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 263.300000 0.600000 263.500000 ;
    END
  END mem_in_core1[31]
  PIN mem_in_core1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 264.100000 0.600000 264.300000 ;
    END
  END mem_in_core1[30]
  PIN mem_in_core1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 264.900000 0.600000 265.100000 ;
    END
  END mem_in_core1[29]
  PIN mem_in_core1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 265.700000 0.600000 265.900000 ;
    END
  END mem_in_core1[28]
  PIN mem_in_core1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 266.500000 0.600000 266.700000 ;
    END
  END mem_in_core1[27]
  PIN mem_in_core1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 267.300000 0.600000 267.500000 ;
    END
  END mem_in_core1[26]
  PIN mem_in_core1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 268.100000 0.600000 268.300000 ;
    END
  END mem_in_core1[25]
  PIN mem_in_core1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 268.900000 0.600000 269.100000 ;
    END
  END mem_in_core1[24]
  PIN mem_in_core1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 269.700000 0.600000 269.900000 ;
    END
  END mem_in_core1[23]
  PIN mem_in_core1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 270.500000 0.600000 270.700000 ;
    END
  END mem_in_core1[22]
  PIN mem_in_core1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 271.300000 0.600000 271.500000 ;
    END
  END mem_in_core1[21]
  PIN mem_in_core1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 272.100000 0.600000 272.300000 ;
    END
  END mem_in_core1[20]
  PIN mem_in_core1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 272.900000 0.600000 273.100000 ;
    END
  END mem_in_core1[19]
  PIN mem_in_core1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 273.700000 0.600000 273.900000 ;
    END
  END mem_in_core1[18]
  PIN mem_in_core1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 274.500000 0.600000 274.700000 ;
    END
  END mem_in_core1[17]
  PIN mem_in_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 275.300000 0.600000 275.500000 ;
    END
  END mem_in_core1[16]
  PIN mem_in_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 276.100000 0.600000 276.300000 ;
    END
  END mem_in_core1[15]
  PIN mem_in_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 276.900000 0.600000 277.100000 ;
    END
  END mem_in_core1[14]
  PIN mem_in_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 277.700000 0.600000 277.900000 ;
    END
  END mem_in_core1[13]
  PIN mem_in_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 278.500000 0.600000 278.700000 ;
    END
  END mem_in_core1[12]
  PIN mem_in_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 279.300000 0.600000 279.500000 ;
    END
  END mem_in_core1[11]
  PIN mem_in_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 280.100000 0.600000 280.300000 ;
    END
  END mem_in_core1[10]
  PIN mem_in_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 280.900000 0.600000 281.100000 ;
    END
  END mem_in_core1[9]
  PIN mem_in_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 281.700000 0.600000 281.900000 ;
    END
  END mem_in_core1[8]
  PIN mem_in_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 282.500000 0.600000 282.700000 ;
    END
  END mem_in_core1[7]
  PIN mem_in_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 283.300000 0.600000 283.500000 ;
    END
  END mem_in_core1[6]
  PIN mem_in_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 284.100000 0.600000 284.300000 ;
    END
  END mem_in_core1[5]
  PIN mem_in_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 284.900000 0.600000 285.100000 ;
    END
  END mem_in_core1[4]
  PIN mem_in_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 285.700000 0.600000 285.900000 ;
    END
  END mem_in_core1[3]
  PIN mem_in_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 286.500000 0.600000 286.700000 ;
    END
  END mem_in_core1[2]
  PIN mem_in_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 287.300000 0.600000 287.500000 ;
    END
  END mem_in_core1[1]
  PIN mem_in_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 288.100000 0.600000 288.300000 ;
    END
  END mem_in_core1[0]
  PIN inst_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 236.100000 0.600000 236.300000 ;
    END
  END inst_core1[16]
  PIN inst_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 236.900000 0.600000 237.100000 ;
    END
  END inst_core1[15]
  PIN inst_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 237.700000 0.600000 237.900000 ;
    END
  END inst_core1[14]
  PIN inst_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 238.500000 0.600000 238.700000 ;
    END
  END inst_core1[13]
  PIN inst_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 239.300000 0.600000 239.500000 ;
    END
  END inst_core1[12]
  PIN inst_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 240.100000 0.600000 240.300000 ;
    END
  END inst_core1[11]
  PIN inst_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 240.900000 0.600000 241.100000 ;
    END
  END inst_core1[10]
  PIN inst_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 241.700000 0.600000 241.900000 ;
    END
  END inst_core1[9]
  PIN inst_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 242.500000 0.600000 242.700000 ;
    END
  END inst_core1[8]
  PIN inst_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 243.300000 0.600000 243.500000 ;
    END
  END inst_core1[7]
  PIN inst_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 244.100000 0.600000 244.300000 ;
    END
  END inst_core1[6]
  PIN inst_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 244.900000 0.600000 245.100000 ;
    END
  END inst_core1[5]
  PIN inst_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 245.700000 0.600000 245.900000 ;
    END
  END inst_core1[4]
  PIN inst_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 246.500000 0.600000 246.700000 ;
    END
  END inst_core1[3]
  PIN inst_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 247.300000 0.600000 247.500000 ;
    END
  END inst_core1[2]
  PIN inst_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 248.100000 0.600000 248.300000 ;
    END
  END inst_core1[1]
  PIN inst_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 248.900000 0.600000 249.100000 ;
    END
  END inst_core1[0]
  PIN out_core1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.000000 0.000000 213.200000 0.600000 ;
    END
  END out_core1[87]
  PIN out_core1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.800000 0.000000 214.000000 0.600000 ;
    END
  END out_core1[86]
  PIN out_core1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.600000 0.000000 214.800000 0.600000 ;
    END
  END out_core1[85]
  PIN out_core1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.400000 0.000000 215.600000 0.600000 ;
    END
  END out_core1[84]
  PIN out_core1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.200000 0.000000 216.400000 0.600000 ;
    END
  END out_core1[83]
  PIN out_core1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.000000 0.000000 217.200000 0.600000 ;
    END
  END out_core1[82]
  PIN out_core1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.800000 0.000000 218.000000 0.600000 ;
    END
  END out_core1[81]
  PIN out_core1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.600000 0.000000 218.800000 0.600000 ;
    END
  END out_core1[80]
  PIN out_core1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.400000 0.000000 219.600000 0.600000 ;
    END
  END out_core1[79]
  PIN out_core1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.200000 0.000000 220.400000 0.600000 ;
    END
  END out_core1[78]
  PIN out_core1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 221.000000 0.000000 221.200000 0.600000 ;
    END
  END out_core1[77]
  PIN out_core1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 221.800000 0.000000 222.000000 0.600000 ;
    END
  END out_core1[76]
  PIN out_core1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.600000 0.000000 222.800000 0.600000 ;
    END
  END out_core1[75]
  PIN out_core1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.400000 0.000000 223.600000 0.600000 ;
    END
  END out_core1[74]
  PIN out_core1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.200000 0.000000 224.400000 0.600000 ;
    END
  END out_core1[73]
  PIN out_core1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 225.000000 0.000000 225.200000 0.600000 ;
    END
  END out_core1[72]
  PIN out_core1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 225.800000 0.000000 226.000000 0.600000 ;
    END
  END out_core1[71]
  PIN out_core1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.600000 0.000000 226.800000 0.600000 ;
    END
  END out_core1[70]
  PIN out_core1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.400000 0.000000 227.600000 0.600000 ;
    END
  END out_core1[69]
  PIN out_core1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.200000 0.000000 228.400000 0.600000 ;
    END
  END out_core1[68]
  PIN out_core1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.000000 0.000000 229.200000 0.600000 ;
    END
  END out_core1[67]
  PIN out_core1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.800000 0.000000 230.000000 0.600000 ;
    END
  END out_core1[66]
  PIN out_core1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.600000 0.000000 230.800000 0.600000 ;
    END
  END out_core1[65]
  PIN out_core1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.400000 0.000000 231.600000 0.600000 ;
    END
  END out_core1[64]
  PIN out_core1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.200000 0.000000 232.400000 0.600000 ;
    END
  END out_core1[63]
  PIN out_core1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.000000 0.000000 233.200000 0.600000 ;
    END
  END out_core1[62]
  PIN out_core1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.800000 0.000000 234.000000 0.600000 ;
    END
  END out_core1[61]
  PIN out_core1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.600000 0.000000 234.800000 0.600000 ;
    END
  END out_core1[60]
  PIN out_core1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.400000 0.000000 235.600000 0.600000 ;
    END
  END out_core1[59]
  PIN out_core1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 236.200000 0.000000 236.400000 0.600000 ;
    END
  END out_core1[58]
  PIN out_core1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.000000 0.000000 237.200000 0.600000 ;
    END
  END out_core1[57]
  PIN out_core1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.800000 0.000000 238.000000 0.600000 ;
    END
  END out_core1[56]
  PIN out_core1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.600000 0.000000 238.800000 0.600000 ;
    END
  END out_core1[55]
  PIN out_core1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 239.400000 0.000000 239.600000 0.600000 ;
    END
  END out_core1[54]
  PIN out_core1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.200000 0.000000 240.400000 0.600000 ;
    END
  END out_core1[53]
  PIN out_core1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.000000 0.000000 241.200000 0.600000 ;
    END
  END out_core1[52]
  PIN out_core1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.800000 0.000000 242.000000 0.600000 ;
    END
  END out_core1[51]
  PIN out_core1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 242.600000 0.000000 242.800000 0.600000 ;
    END
  END out_core1[50]
  PIN out_core1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.400000 0.000000 243.600000 0.600000 ;
    END
  END out_core1[49]
  PIN out_core1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.200000 0.000000 244.400000 0.600000 ;
    END
  END out_core1[48]
  PIN out_core1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.000000 0.000000 245.200000 0.600000 ;
    END
  END out_core1[47]
  PIN out_core1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.800000 0.000000 246.000000 0.600000 ;
    END
  END out_core1[46]
  PIN out_core1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.600000 0.000000 246.800000 0.600000 ;
    END
  END out_core1[45]
  PIN out_core1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.400000 0.000000 247.600000 0.600000 ;
    END
  END out_core1[44]
  PIN out_core1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.200000 0.000000 248.400000 0.600000 ;
    END
  END out_core1[43]
  PIN out_core1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 249.000000 0.000000 249.200000 0.600000 ;
    END
  END out_core1[42]
  PIN out_core1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 249.800000 0.000000 250.000000 0.600000 ;
    END
  END out_core1[41]
  PIN out_core1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.600000 0.000000 250.800000 0.600000 ;
    END
  END out_core1[40]
  PIN out_core1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.400000 0.000000 251.600000 0.600000 ;
    END
  END out_core1[39]
  PIN out_core1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.200000 0.000000 252.400000 0.600000 ;
    END
  END out_core1[38]
  PIN out_core1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 253.000000 0.000000 253.200000 0.600000 ;
    END
  END out_core1[37]
  PIN out_core1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 253.800000 0.000000 254.000000 0.600000 ;
    END
  END out_core1[36]
  PIN out_core1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 254.600000 0.000000 254.800000 0.600000 ;
    END
  END out_core1[35]
  PIN out_core1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.400000 0.000000 255.600000 0.600000 ;
    END
  END out_core1[34]
  PIN out_core1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.200000 0.000000 256.400000 0.600000 ;
    END
  END out_core1[33]
  PIN out_core1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 257.000000 0.000000 257.200000 0.600000 ;
    END
  END out_core1[32]
  PIN out_core1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 257.800000 0.000000 258.000000 0.600000 ;
    END
  END out_core1[31]
  PIN out_core1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.600000 0.000000 258.800000 0.600000 ;
    END
  END out_core1[30]
  PIN out_core1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.400000 0.000000 259.600000 0.600000 ;
    END
  END out_core1[29]
  PIN out_core1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.200000 0.000000 260.400000 0.600000 ;
    END
  END out_core1[28]
  PIN out_core1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.000000 0.000000 261.200000 0.600000 ;
    END
  END out_core1[27]
  PIN out_core1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.800000 0.000000 262.000000 0.600000 ;
    END
  END out_core1[26]
  PIN out_core1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.600000 0.000000 262.800000 0.600000 ;
    END
  END out_core1[25]
  PIN out_core1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.400000 0.000000 263.600000 0.600000 ;
    END
  END out_core1[24]
  PIN out_core1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 264.200000 0.000000 264.400000 0.600000 ;
    END
  END out_core1[23]
  PIN out_core1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.000000 0.000000 265.200000 0.600000 ;
    END
  END out_core1[22]
  PIN out_core1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.800000 0.000000 266.000000 0.600000 ;
    END
  END out_core1[21]
  PIN out_core1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 266.600000 0.000000 266.800000 0.600000 ;
    END
  END out_core1[20]
  PIN out_core1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.400000 0.000000 267.600000 0.600000 ;
    END
  END out_core1[19]
  PIN out_core1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.200000 0.000000 268.400000 0.600000 ;
    END
  END out_core1[18]
  PIN out_core1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 269.000000 0.000000 269.200000 0.600000 ;
    END
  END out_core1[17]
  PIN out_core1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 269.800000 0.000000 270.000000 0.600000 ;
    END
  END out_core1[16]
  PIN out_core1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.600000 0.000000 270.800000 0.600000 ;
    END
  END out_core1[15]
  PIN out_core1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.400000 0.000000 271.600000 0.600000 ;
    END
  END out_core1[14]
  PIN out_core1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 272.200000 0.000000 272.400000 0.600000 ;
    END
  END out_core1[13]
  PIN out_core1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.000000 0.000000 273.200000 0.600000 ;
    END
  END out_core1[12]
  PIN out_core1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.800000 0.000000 274.000000 0.600000 ;
    END
  END out_core1[11]
  PIN out_core1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.600000 0.000000 274.800000 0.600000 ;
    END
  END out_core1[10]
  PIN out_core1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.400000 0.000000 275.600000 0.600000 ;
    END
  END out_core1[9]
  PIN out_core1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 276.200000 0.000000 276.400000 0.600000 ;
    END
  END out_core1[8]
  PIN out_core1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.000000 0.000000 277.200000 0.600000 ;
    END
  END out_core1[7]
  PIN out_core1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.800000 0.000000 278.000000 0.600000 ;
    END
  END out_core1[6]
  PIN out_core1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.600000 0.000000 278.800000 0.600000 ;
    END
  END out_core1[5]
  PIN out_core1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.400000 0.000000 279.600000 0.600000 ;
    END
  END out_core1[4]
  PIN out_core1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.200000 0.000000 280.400000 0.600000 ;
    END
  END out_core1[3]
  PIN out_core1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.000000 0.000000 281.200000 0.600000 ;
    END
  END out_core1[2]
  PIN out_core1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.800000 0.000000 282.000000 0.600000 ;
    END
  END out_core1[1]
  PIN out_core1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.600000 0.000000 282.800000 0.600000 ;
    END
  END out_core1[0]
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 232.100000 0.600000 232.300000 ;
    END
  END clk2
  PIN rst2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 235.300000 0.600000 235.500000 ;
    END
  END rst2
  PIN mem_in_core2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 288.900000 0.600000 289.100000 ;
    END
  END mem_in_core2[31]
  PIN mem_in_core2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 289.700000 0.600000 289.900000 ;
    END
  END mem_in_core2[30]
  PIN mem_in_core2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 290.500000 0.600000 290.700000 ;
    END
  END mem_in_core2[29]
  PIN mem_in_core2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 291.300000 0.600000 291.500000 ;
    END
  END mem_in_core2[28]
  PIN mem_in_core2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 292.100000 0.600000 292.300000 ;
    END
  END mem_in_core2[27]
  PIN mem_in_core2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 292.900000 0.600000 293.100000 ;
    END
  END mem_in_core2[26]
  PIN mem_in_core2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 293.700000 0.600000 293.900000 ;
    END
  END mem_in_core2[25]
  PIN mem_in_core2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 294.500000 0.600000 294.700000 ;
    END
  END mem_in_core2[24]
  PIN mem_in_core2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 295.300000 0.600000 295.500000 ;
    END
  END mem_in_core2[23]
  PIN mem_in_core2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 296.100000 0.600000 296.300000 ;
    END
  END mem_in_core2[22]
  PIN mem_in_core2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 296.900000 0.600000 297.100000 ;
    END
  END mem_in_core2[21]
  PIN mem_in_core2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 297.700000 0.600000 297.900000 ;
    END
  END mem_in_core2[20]
  PIN mem_in_core2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 298.500000 0.600000 298.700000 ;
    END
  END mem_in_core2[19]
  PIN mem_in_core2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 299.300000 0.600000 299.500000 ;
    END
  END mem_in_core2[18]
  PIN mem_in_core2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 300.100000 0.600000 300.300000 ;
    END
  END mem_in_core2[17]
  PIN mem_in_core2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 300.900000 0.600000 301.100000 ;
    END
  END mem_in_core2[16]
  PIN mem_in_core2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 301.700000 0.600000 301.900000 ;
    END
  END mem_in_core2[15]
  PIN mem_in_core2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 302.500000 0.600000 302.700000 ;
    END
  END mem_in_core2[14]
  PIN mem_in_core2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 303.300000 0.600000 303.500000 ;
    END
  END mem_in_core2[13]
  PIN mem_in_core2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.100000 0.600000 304.300000 ;
    END
  END mem_in_core2[12]
  PIN mem_in_core2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.900000 0.600000 305.100000 ;
    END
  END mem_in_core2[11]
  PIN mem_in_core2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 305.700000 0.600000 305.900000 ;
    END
  END mem_in_core2[10]
  PIN mem_in_core2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 306.500000 0.600000 306.700000 ;
    END
  END mem_in_core2[9]
  PIN mem_in_core2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 307.300000 0.600000 307.500000 ;
    END
  END mem_in_core2[8]
  PIN mem_in_core2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 308.100000 0.600000 308.300000 ;
    END
  END mem_in_core2[7]
  PIN mem_in_core2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 308.900000 0.600000 309.100000 ;
    END
  END mem_in_core2[6]
  PIN mem_in_core2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 309.700000 0.600000 309.900000 ;
    END
  END mem_in_core2[5]
  PIN mem_in_core2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 310.500000 0.600000 310.700000 ;
    END
  END mem_in_core2[4]
  PIN mem_in_core2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 311.300000 0.600000 311.500000 ;
    END
  END mem_in_core2[3]
  PIN mem_in_core2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 312.100000 0.600000 312.300000 ;
    END
  END mem_in_core2[2]
  PIN mem_in_core2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 312.900000 0.600000 313.100000 ;
    END
  END mem_in_core2[1]
  PIN mem_in_core2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 313.700000 0.600000 313.900000 ;
    END
  END mem_in_core2[0]
  PIN inst_core2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 249.700000 0.600000 249.900000 ;
    END
  END inst_core2[16]
  PIN inst_core2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 250.500000 0.600000 250.700000 ;
    END
  END inst_core2[15]
  PIN inst_core2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 251.300000 0.600000 251.500000 ;
    END
  END inst_core2[14]
  PIN inst_core2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 252.100000 0.600000 252.300000 ;
    END
  END inst_core2[13]
  PIN inst_core2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 252.900000 0.600000 253.100000 ;
    END
  END inst_core2[12]
  PIN inst_core2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 253.700000 0.600000 253.900000 ;
    END
  END inst_core2[11]
  PIN inst_core2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 254.500000 0.600000 254.700000 ;
    END
  END inst_core2[10]
  PIN inst_core2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 255.300000 0.600000 255.500000 ;
    END
  END inst_core2[9]
  PIN inst_core2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 256.100000 0.600000 256.300000 ;
    END
  END inst_core2[8]
  PIN inst_core2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 256.900000 0.600000 257.100000 ;
    END
  END inst_core2[7]
  PIN inst_core2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 257.700000 0.600000 257.900000 ;
    END
  END inst_core2[6]
  PIN inst_core2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 258.500000 0.600000 258.700000 ;
    END
  END inst_core2[5]
  PIN inst_core2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 259.300000 0.600000 259.500000 ;
    END
  END inst_core2[4]
  PIN inst_core2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 260.100000 0.600000 260.300000 ;
    END
  END inst_core2[3]
  PIN inst_core2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 260.900000 0.600000 261.100000 ;
    END
  END inst_core2[2]
  PIN inst_core2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 261.700000 0.600000 261.900000 ;
    END
  END inst_core2[1]
  PIN inst_core2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 262.500000 0.600000 262.700000 ;
    END
  END inst_core2[0]
  PIN out_core2[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.400000 0.000000 283.600000 0.600000 ;
    END
  END out_core2[87]
  PIN out_core2[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284.200000 0.000000 284.400000 0.600000 ;
    END
  END out_core2[86]
  PIN out_core2[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.000000 0.000000 285.200000 0.600000 ;
    END
  END out_core2[85]
  PIN out_core2[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.800000 0.000000 286.000000 0.600000 ;
    END
  END out_core2[84]
  PIN out_core2[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 286.600000 0.000000 286.800000 0.600000 ;
    END
  END out_core2[83]
  PIN out_core2[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.400000 0.000000 287.600000 0.600000 ;
    END
  END out_core2[82]
  PIN out_core2[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.200000 0.000000 288.400000 0.600000 ;
    END
  END out_core2[81]
  PIN out_core2[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.000000 0.000000 289.200000 0.600000 ;
    END
  END out_core2[80]
  PIN out_core2[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.800000 0.000000 290.000000 0.600000 ;
    END
  END out_core2[79]
  PIN out_core2[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 290.600000 0.000000 290.800000 0.600000 ;
    END
  END out_core2[78]
  PIN out_core2[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.400000 0.000000 291.600000 0.600000 ;
    END
  END out_core2[77]
  PIN out_core2[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 292.200000 0.000000 292.400000 0.600000 ;
    END
  END out_core2[76]
  PIN out_core2[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 293.000000 0.000000 293.200000 0.600000 ;
    END
  END out_core2[75]
  PIN out_core2[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 293.800000 0.000000 294.000000 0.600000 ;
    END
  END out_core2[74]
  PIN out_core2[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 294.600000 0.000000 294.800000 0.600000 ;
    END
  END out_core2[73]
  PIN out_core2[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.400000 0.000000 295.600000 0.600000 ;
    END
  END out_core2[72]
  PIN out_core2[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 296.200000 0.000000 296.400000 0.600000 ;
    END
  END out_core2[71]
  PIN out_core2[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.000000 0.000000 297.200000 0.600000 ;
    END
  END out_core2[70]
  PIN out_core2[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.800000 0.000000 298.000000 0.600000 ;
    END
  END out_core2[69]
  PIN out_core2[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 298.600000 0.000000 298.800000 0.600000 ;
    END
  END out_core2[68]
  PIN out_core2[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.400000 0.000000 299.600000 0.600000 ;
    END
  END out_core2[67]
  PIN out_core2[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.200000 0.000000 300.400000 0.600000 ;
    END
  END out_core2[66]
  PIN out_core2[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 301.000000 0.000000 301.200000 0.600000 ;
    END
  END out_core2[65]
  PIN out_core2[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 301.800000 0.000000 302.000000 0.600000 ;
    END
  END out_core2[64]
  PIN out_core2[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.600000 0.000000 302.800000 0.600000 ;
    END
  END out_core2[63]
  PIN out_core2[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.400000 0.000000 303.600000 0.600000 ;
    END
  END out_core2[62]
  PIN out_core2[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 304.200000 0.000000 304.400000 0.600000 ;
    END
  END out_core2[61]
  PIN out_core2[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.000000 0.000000 305.200000 0.600000 ;
    END
  END out_core2[60]
  PIN out_core2[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.800000 0.000000 306.000000 0.600000 ;
    END
  END out_core2[59]
  PIN out_core2[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.600000 0.000000 306.800000 0.600000 ;
    END
  END out_core2[58]
  PIN out_core2[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.400000 0.000000 307.600000 0.600000 ;
    END
  END out_core2[57]
  PIN out_core2[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.200000 0.000000 308.400000 0.600000 ;
    END
  END out_core2[56]
  PIN out_core2[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.000000 0.000000 309.200000 0.600000 ;
    END
  END out_core2[55]
  PIN out_core2[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.800000 0.000000 310.000000 0.600000 ;
    END
  END out_core2[54]
  PIN out_core2[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.600000 0.000000 310.800000 0.600000 ;
    END
  END out_core2[53]
  PIN out_core2[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.400000 0.000000 311.600000 0.600000 ;
    END
  END out_core2[52]
  PIN out_core2[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.200000 0.000000 312.400000 0.600000 ;
    END
  END out_core2[51]
  PIN out_core2[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.000000 0.000000 313.200000 0.600000 ;
    END
  END out_core2[50]
  PIN out_core2[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.800000 0.000000 314.000000 0.600000 ;
    END
  END out_core2[49]
  PIN out_core2[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.600000 0.000000 314.800000 0.600000 ;
    END
  END out_core2[48]
  PIN out_core2[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.400000 0.000000 315.600000 0.600000 ;
    END
  END out_core2[47]
  PIN out_core2[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.200000 0.000000 316.400000 0.600000 ;
    END
  END out_core2[46]
  PIN out_core2[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.000000 0.000000 317.200000 0.600000 ;
    END
  END out_core2[45]
  PIN out_core2[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.800000 0.000000 318.000000 0.600000 ;
    END
  END out_core2[44]
  PIN out_core2[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.600000 0.000000 318.800000 0.600000 ;
    END
  END out_core2[43]
  PIN out_core2[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.400000 0.000000 319.600000 0.600000 ;
    END
  END out_core2[42]
  PIN out_core2[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.200000 0.000000 320.400000 0.600000 ;
    END
  END out_core2[41]
  PIN out_core2[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.000000 0.000000 321.200000 0.600000 ;
    END
  END out_core2[40]
  PIN out_core2[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.800000 0.000000 322.000000 0.600000 ;
    END
  END out_core2[39]
  PIN out_core2[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.600000 0.000000 322.800000 0.600000 ;
    END
  END out_core2[38]
  PIN out_core2[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.400000 0.000000 323.600000 0.600000 ;
    END
  END out_core2[37]
  PIN out_core2[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.200000 0.000000 324.400000 0.600000 ;
    END
  END out_core2[36]
  PIN out_core2[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.000000 0.000000 325.200000 0.600000 ;
    END
  END out_core2[35]
  PIN out_core2[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.800000 0.000000 326.000000 0.600000 ;
    END
  END out_core2[34]
  PIN out_core2[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.600000 0.000000 326.800000 0.600000 ;
    END
  END out_core2[33]
  PIN out_core2[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.400000 0.000000 327.600000 0.600000 ;
    END
  END out_core2[32]
  PIN out_core2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.200000 0.000000 328.400000 0.600000 ;
    END
  END out_core2[31]
  PIN out_core2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.000000 0.000000 329.200000 0.600000 ;
    END
  END out_core2[30]
  PIN out_core2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.800000 0.000000 330.000000 0.600000 ;
    END
  END out_core2[29]
  PIN out_core2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.600000 0.000000 330.800000 0.600000 ;
    END
  END out_core2[28]
  PIN out_core2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.400000 0.000000 331.600000 0.600000 ;
    END
  END out_core2[27]
  PIN out_core2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.200000 0.000000 332.400000 0.600000 ;
    END
  END out_core2[26]
  PIN out_core2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.000000 0.000000 333.200000 0.600000 ;
    END
  END out_core2[25]
  PIN out_core2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.800000 0.000000 334.000000 0.600000 ;
    END
  END out_core2[24]
  PIN out_core2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.600000 0.000000 334.800000 0.600000 ;
    END
  END out_core2[23]
  PIN out_core2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.400000 0.000000 335.600000 0.600000 ;
    END
  END out_core2[22]
  PIN out_core2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.200000 0.000000 336.400000 0.600000 ;
    END
  END out_core2[21]
  PIN out_core2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.000000 0.000000 337.200000 0.600000 ;
    END
  END out_core2[20]
  PIN out_core2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.800000 0.000000 338.000000 0.600000 ;
    END
  END out_core2[19]
  PIN out_core2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.600000 0.000000 338.800000 0.600000 ;
    END
  END out_core2[18]
  PIN out_core2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.400000 0.000000 339.600000 0.600000 ;
    END
  END out_core2[17]
  PIN out_core2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.200000 0.000000 340.400000 0.600000 ;
    END
  END out_core2[16]
  PIN out_core2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.000000 0.000000 341.200000 0.600000 ;
    END
  END out_core2[15]
  PIN out_core2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.800000 0.000000 342.000000 0.600000 ;
    END
  END out_core2[14]
  PIN out_core2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.600000 0.000000 342.800000 0.600000 ;
    END
  END out_core2[13]
  PIN out_core2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.400000 0.000000 343.600000 0.600000 ;
    END
  END out_core2[12]
  PIN out_core2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.200000 0.000000 344.400000 0.600000 ;
    END
  END out_core2[11]
  PIN out_core2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.000000 0.000000 345.200000 0.600000 ;
    END
  END out_core2[10]
  PIN out_core2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.800000 0.000000 346.000000 0.600000 ;
    END
  END out_core2[9]
  PIN out_core2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.600000 0.000000 346.800000 0.600000 ;
    END
  END out_core2[8]
  PIN out_core2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.400000 0.000000 347.600000 0.600000 ;
    END
  END out_core2[7]
  PIN out_core2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.200000 0.000000 348.400000 0.600000 ;
    END
  END out_core2[6]
  PIN out_core2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.000000 0.000000 349.200000 0.600000 ;
    END
  END out_core2[5]
  PIN out_core2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.800000 0.000000 350.000000 0.600000 ;
    END
  END out_core2[4]
  PIN out_core2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.600000 0.000000 350.800000 0.600000 ;
    END
  END out_core2[3]
  PIN out_core2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.400000 0.000000 351.600000 0.600000 ;
    END
  END out_core2[2]
  PIN out_core2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.200000 0.000000 352.400000 0.600000 ;
    END
  END out_core2[1]
  PIN out_core2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.000000 0.000000 353.200000 0.600000 ;
    END
  END out_core2[0]
  PIN core_gate1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 232.900000 0.600000 233.100000 ;
    END
  END core_gate1
  PIN core_gate2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 233.700000 0.600000 233.900000 ;
    END
  END core_gate2
  PIN s_valid1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.000000 0.000000 193.200000 0.600000 ;
    END
  END s_valid1
  PIN s_valid2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.800000 0.000000 194.000000 0.600000 ;
    END
  END s_valid2
  PIN psum_norm_1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.400000 0.000000 195.600000 0.600000 ;
    END
  END psum_norm_1[10]
  PIN psum_norm_1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.200000 0.000000 196.400000 0.600000 ;
    END
  END psum_norm_1[9]
  PIN psum_norm_1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.000000 0.000000 197.200000 0.600000 ;
    END
  END psum_norm_1[8]
  PIN psum_norm_1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.800000 0.000000 198.000000 0.600000 ;
    END
  END psum_norm_1[7]
  PIN psum_norm_1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.600000 0.000000 198.800000 0.600000 ;
    END
  END psum_norm_1[6]
  PIN psum_norm_1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.400000 0.000000 199.600000 0.600000 ;
    END
  END psum_norm_1[5]
  PIN psum_norm_1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.200000 0.000000 200.400000 0.600000 ;
    END
  END psum_norm_1[4]
  PIN psum_norm_1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.000000 0.000000 201.200000 0.600000 ;
    END
  END psum_norm_1[3]
  PIN psum_norm_1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.800000 0.000000 202.000000 0.600000 ;
    END
  END psum_norm_1[2]
  PIN psum_norm_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.600000 0.000000 202.800000 0.600000 ;
    END
  END psum_norm_1[1]
  PIN psum_norm_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.400000 0.000000 203.600000 0.600000 ;
    END
  END psum_norm_1[0]
  PIN psum_norm_2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.200000 0.000000 204.400000 0.600000 ;
    END
  END psum_norm_2[10]
  PIN psum_norm_2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.000000 0.000000 205.200000 0.600000 ;
    END
  END psum_norm_2[9]
  PIN psum_norm_2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.800000 0.000000 206.000000 0.600000 ;
    END
  END psum_norm_2[8]
  PIN psum_norm_2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.600000 0.000000 206.800000 0.600000 ;
    END
  END psum_norm_2[7]
  PIN psum_norm_2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.400000 0.000000 207.600000 0.600000 ;
    END
  END psum_norm_2[6]
  PIN psum_norm_2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.200000 0.000000 208.400000 0.600000 ;
    END
  END psum_norm_2[5]
  PIN psum_norm_2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.000000 0.000000 209.200000 0.600000 ;
    END
  END psum_norm_2[4]
  PIN psum_norm_2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.800000 0.000000 210.000000 0.600000 ;
    END
  END psum_norm_2[3]
  PIN psum_norm_2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.600000 0.000000 210.800000 0.600000 ;
    END
  END psum_norm_2[2]
  PIN psum_norm_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.400000 0.000000 211.600000 0.600000 ;
    END
  END psum_norm_2[1]
  PIN psum_norm_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.200000 0.000000 212.400000 0.600000 ;
    END
  END psum_norm_2[0]
  PIN norm_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.600000 0.000000 194.800000 0.600000 ;
    END
  END norm_valid
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 546.600000 545.600000 ;
    LAYER M2 ;
      RECT 0.000000 0.700000 546.600000 545.600000 ;
      RECT 353.300000 0.000000 546.600000 0.700000 ;
      RECT 352.500000 0.000000 352.900000 0.700000 ;
      RECT 351.700000 0.000000 352.100000 0.700000 ;
      RECT 350.900000 0.000000 351.300000 0.700000 ;
      RECT 350.100000 0.000000 350.500000 0.700000 ;
      RECT 349.300000 0.000000 349.700000 0.700000 ;
      RECT 348.500000 0.000000 348.900000 0.700000 ;
      RECT 347.700000 0.000000 348.100000 0.700000 ;
      RECT 346.900000 0.000000 347.300000 0.700000 ;
      RECT 346.100000 0.000000 346.500000 0.700000 ;
      RECT 345.300000 0.000000 345.700000 0.700000 ;
      RECT 344.500000 0.000000 344.900000 0.700000 ;
      RECT 343.700000 0.000000 344.100000 0.700000 ;
      RECT 342.900000 0.000000 343.300000 0.700000 ;
      RECT 342.100000 0.000000 342.500000 0.700000 ;
      RECT 341.300000 0.000000 341.700000 0.700000 ;
      RECT 340.500000 0.000000 340.900000 0.700000 ;
      RECT 339.700000 0.000000 340.100000 0.700000 ;
      RECT 338.900000 0.000000 339.300000 0.700000 ;
      RECT 338.100000 0.000000 338.500000 0.700000 ;
      RECT 337.300000 0.000000 337.700000 0.700000 ;
      RECT 336.500000 0.000000 336.900000 0.700000 ;
      RECT 335.700000 0.000000 336.100000 0.700000 ;
      RECT 334.900000 0.000000 335.300000 0.700000 ;
      RECT 334.100000 0.000000 334.500000 0.700000 ;
      RECT 333.300000 0.000000 333.700000 0.700000 ;
      RECT 332.500000 0.000000 332.900000 0.700000 ;
      RECT 331.700000 0.000000 332.100000 0.700000 ;
      RECT 330.900000 0.000000 331.300000 0.700000 ;
      RECT 330.100000 0.000000 330.500000 0.700000 ;
      RECT 329.300000 0.000000 329.700000 0.700000 ;
      RECT 328.500000 0.000000 328.900000 0.700000 ;
      RECT 327.700000 0.000000 328.100000 0.700000 ;
      RECT 326.900000 0.000000 327.300000 0.700000 ;
      RECT 326.100000 0.000000 326.500000 0.700000 ;
      RECT 325.300000 0.000000 325.700000 0.700000 ;
      RECT 324.500000 0.000000 324.900000 0.700000 ;
      RECT 323.700000 0.000000 324.100000 0.700000 ;
      RECT 322.900000 0.000000 323.300000 0.700000 ;
      RECT 322.100000 0.000000 322.500000 0.700000 ;
      RECT 321.300000 0.000000 321.700000 0.700000 ;
      RECT 320.500000 0.000000 320.900000 0.700000 ;
      RECT 319.700000 0.000000 320.100000 0.700000 ;
      RECT 318.900000 0.000000 319.300000 0.700000 ;
      RECT 318.100000 0.000000 318.500000 0.700000 ;
      RECT 317.300000 0.000000 317.700000 0.700000 ;
      RECT 316.500000 0.000000 316.900000 0.700000 ;
      RECT 315.700000 0.000000 316.100000 0.700000 ;
      RECT 314.900000 0.000000 315.300000 0.700000 ;
      RECT 314.100000 0.000000 314.500000 0.700000 ;
      RECT 313.300000 0.000000 313.700000 0.700000 ;
      RECT 312.500000 0.000000 312.900000 0.700000 ;
      RECT 311.700000 0.000000 312.100000 0.700000 ;
      RECT 310.900000 0.000000 311.300000 0.700000 ;
      RECT 310.100000 0.000000 310.500000 0.700000 ;
      RECT 309.300000 0.000000 309.700000 0.700000 ;
      RECT 308.500000 0.000000 308.900000 0.700000 ;
      RECT 307.700000 0.000000 308.100000 0.700000 ;
      RECT 306.900000 0.000000 307.300000 0.700000 ;
      RECT 306.100000 0.000000 306.500000 0.700000 ;
      RECT 305.300000 0.000000 305.700000 0.700000 ;
      RECT 304.500000 0.000000 304.900000 0.700000 ;
      RECT 303.700000 0.000000 304.100000 0.700000 ;
      RECT 302.900000 0.000000 303.300000 0.700000 ;
      RECT 302.100000 0.000000 302.500000 0.700000 ;
      RECT 301.300000 0.000000 301.700000 0.700000 ;
      RECT 300.500000 0.000000 300.900000 0.700000 ;
      RECT 299.700000 0.000000 300.100000 0.700000 ;
      RECT 298.900000 0.000000 299.300000 0.700000 ;
      RECT 298.100000 0.000000 298.500000 0.700000 ;
      RECT 297.300000 0.000000 297.700000 0.700000 ;
      RECT 296.500000 0.000000 296.900000 0.700000 ;
      RECT 295.700000 0.000000 296.100000 0.700000 ;
      RECT 294.900000 0.000000 295.300000 0.700000 ;
      RECT 294.100000 0.000000 294.500000 0.700000 ;
      RECT 293.300000 0.000000 293.700000 0.700000 ;
      RECT 292.500000 0.000000 292.900000 0.700000 ;
      RECT 291.700000 0.000000 292.100000 0.700000 ;
      RECT 290.900000 0.000000 291.300000 0.700000 ;
      RECT 290.100000 0.000000 290.500000 0.700000 ;
      RECT 289.300000 0.000000 289.700000 0.700000 ;
      RECT 288.500000 0.000000 288.900000 0.700000 ;
      RECT 287.700000 0.000000 288.100000 0.700000 ;
      RECT 286.900000 0.000000 287.300000 0.700000 ;
      RECT 286.100000 0.000000 286.500000 0.700000 ;
      RECT 285.300000 0.000000 285.700000 0.700000 ;
      RECT 284.500000 0.000000 284.900000 0.700000 ;
      RECT 283.700000 0.000000 284.100000 0.700000 ;
      RECT 282.900000 0.000000 283.300000 0.700000 ;
      RECT 282.100000 0.000000 282.500000 0.700000 ;
      RECT 281.300000 0.000000 281.700000 0.700000 ;
      RECT 280.500000 0.000000 280.900000 0.700000 ;
      RECT 279.700000 0.000000 280.100000 0.700000 ;
      RECT 278.900000 0.000000 279.300000 0.700000 ;
      RECT 278.100000 0.000000 278.500000 0.700000 ;
      RECT 277.300000 0.000000 277.700000 0.700000 ;
      RECT 276.500000 0.000000 276.900000 0.700000 ;
      RECT 275.700000 0.000000 276.100000 0.700000 ;
      RECT 274.900000 0.000000 275.300000 0.700000 ;
      RECT 274.100000 0.000000 274.500000 0.700000 ;
      RECT 273.300000 0.000000 273.700000 0.700000 ;
      RECT 272.500000 0.000000 272.900000 0.700000 ;
      RECT 271.700000 0.000000 272.100000 0.700000 ;
      RECT 270.900000 0.000000 271.300000 0.700000 ;
      RECT 270.100000 0.000000 270.500000 0.700000 ;
      RECT 269.300000 0.000000 269.700000 0.700000 ;
      RECT 268.500000 0.000000 268.900000 0.700000 ;
      RECT 267.700000 0.000000 268.100000 0.700000 ;
      RECT 266.900000 0.000000 267.300000 0.700000 ;
      RECT 266.100000 0.000000 266.500000 0.700000 ;
      RECT 265.300000 0.000000 265.700000 0.700000 ;
      RECT 264.500000 0.000000 264.900000 0.700000 ;
      RECT 263.700000 0.000000 264.100000 0.700000 ;
      RECT 262.900000 0.000000 263.300000 0.700000 ;
      RECT 262.100000 0.000000 262.500000 0.700000 ;
      RECT 261.300000 0.000000 261.700000 0.700000 ;
      RECT 260.500000 0.000000 260.900000 0.700000 ;
      RECT 259.700000 0.000000 260.100000 0.700000 ;
      RECT 258.900000 0.000000 259.300000 0.700000 ;
      RECT 258.100000 0.000000 258.500000 0.700000 ;
      RECT 257.300000 0.000000 257.700000 0.700000 ;
      RECT 256.500000 0.000000 256.900000 0.700000 ;
      RECT 255.700000 0.000000 256.100000 0.700000 ;
      RECT 254.900000 0.000000 255.300000 0.700000 ;
      RECT 254.100000 0.000000 254.500000 0.700000 ;
      RECT 253.300000 0.000000 253.700000 0.700000 ;
      RECT 252.500000 0.000000 252.900000 0.700000 ;
      RECT 251.700000 0.000000 252.100000 0.700000 ;
      RECT 250.900000 0.000000 251.300000 0.700000 ;
      RECT 250.100000 0.000000 250.500000 0.700000 ;
      RECT 249.300000 0.000000 249.700000 0.700000 ;
      RECT 248.500000 0.000000 248.900000 0.700000 ;
      RECT 247.700000 0.000000 248.100000 0.700000 ;
      RECT 246.900000 0.000000 247.300000 0.700000 ;
      RECT 246.100000 0.000000 246.500000 0.700000 ;
      RECT 245.300000 0.000000 245.700000 0.700000 ;
      RECT 244.500000 0.000000 244.900000 0.700000 ;
      RECT 243.700000 0.000000 244.100000 0.700000 ;
      RECT 242.900000 0.000000 243.300000 0.700000 ;
      RECT 242.100000 0.000000 242.500000 0.700000 ;
      RECT 241.300000 0.000000 241.700000 0.700000 ;
      RECT 240.500000 0.000000 240.900000 0.700000 ;
      RECT 239.700000 0.000000 240.100000 0.700000 ;
      RECT 238.900000 0.000000 239.300000 0.700000 ;
      RECT 238.100000 0.000000 238.500000 0.700000 ;
      RECT 237.300000 0.000000 237.700000 0.700000 ;
      RECT 236.500000 0.000000 236.900000 0.700000 ;
      RECT 235.700000 0.000000 236.100000 0.700000 ;
      RECT 234.900000 0.000000 235.300000 0.700000 ;
      RECT 234.100000 0.000000 234.500000 0.700000 ;
      RECT 233.300000 0.000000 233.700000 0.700000 ;
      RECT 232.500000 0.000000 232.900000 0.700000 ;
      RECT 231.700000 0.000000 232.100000 0.700000 ;
      RECT 230.900000 0.000000 231.300000 0.700000 ;
      RECT 230.100000 0.000000 230.500000 0.700000 ;
      RECT 229.300000 0.000000 229.700000 0.700000 ;
      RECT 228.500000 0.000000 228.900000 0.700000 ;
      RECT 227.700000 0.000000 228.100000 0.700000 ;
      RECT 226.900000 0.000000 227.300000 0.700000 ;
      RECT 226.100000 0.000000 226.500000 0.700000 ;
      RECT 225.300000 0.000000 225.700000 0.700000 ;
      RECT 224.500000 0.000000 224.900000 0.700000 ;
      RECT 223.700000 0.000000 224.100000 0.700000 ;
      RECT 222.900000 0.000000 223.300000 0.700000 ;
      RECT 222.100000 0.000000 222.500000 0.700000 ;
      RECT 221.300000 0.000000 221.700000 0.700000 ;
      RECT 220.500000 0.000000 220.900000 0.700000 ;
      RECT 219.700000 0.000000 220.100000 0.700000 ;
      RECT 218.900000 0.000000 219.300000 0.700000 ;
      RECT 218.100000 0.000000 218.500000 0.700000 ;
      RECT 217.300000 0.000000 217.700000 0.700000 ;
      RECT 216.500000 0.000000 216.900000 0.700000 ;
      RECT 215.700000 0.000000 216.100000 0.700000 ;
      RECT 214.900000 0.000000 215.300000 0.700000 ;
      RECT 214.100000 0.000000 214.500000 0.700000 ;
      RECT 213.300000 0.000000 213.700000 0.700000 ;
      RECT 212.500000 0.000000 212.900000 0.700000 ;
      RECT 211.700000 0.000000 212.100000 0.700000 ;
      RECT 210.900000 0.000000 211.300000 0.700000 ;
      RECT 210.100000 0.000000 210.500000 0.700000 ;
      RECT 209.300000 0.000000 209.700000 0.700000 ;
      RECT 208.500000 0.000000 208.900000 0.700000 ;
      RECT 207.700000 0.000000 208.100000 0.700000 ;
      RECT 206.900000 0.000000 207.300000 0.700000 ;
      RECT 206.100000 0.000000 206.500000 0.700000 ;
      RECT 205.300000 0.000000 205.700000 0.700000 ;
      RECT 204.500000 0.000000 204.900000 0.700000 ;
      RECT 203.700000 0.000000 204.100000 0.700000 ;
      RECT 202.900000 0.000000 203.300000 0.700000 ;
      RECT 202.100000 0.000000 202.500000 0.700000 ;
      RECT 201.300000 0.000000 201.700000 0.700000 ;
      RECT 200.500000 0.000000 200.900000 0.700000 ;
      RECT 199.700000 0.000000 200.100000 0.700000 ;
      RECT 198.900000 0.000000 199.300000 0.700000 ;
      RECT 198.100000 0.000000 198.500000 0.700000 ;
      RECT 197.300000 0.000000 197.700000 0.700000 ;
      RECT 196.500000 0.000000 196.900000 0.700000 ;
      RECT 195.700000 0.000000 196.100000 0.700000 ;
      RECT 194.900000 0.000000 195.300000 0.700000 ;
      RECT 194.100000 0.000000 194.500000 0.700000 ;
      RECT 193.300000 0.000000 193.700000 0.700000 ;
      RECT 0.000000 0.000000 192.900000 0.700000 ;
    LAYER M3 ;
      RECT 0.000000 314.000000 546.600000 545.600000 ;
      RECT 0.700000 313.600000 546.600000 314.000000 ;
      RECT 0.000000 313.200000 546.600000 313.600000 ;
      RECT 0.700000 312.800000 546.600000 313.200000 ;
      RECT 0.000000 312.400000 546.600000 312.800000 ;
      RECT 0.700000 312.000000 546.600000 312.400000 ;
      RECT 0.000000 311.600000 546.600000 312.000000 ;
      RECT 0.700000 311.200000 546.600000 311.600000 ;
      RECT 0.000000 310.800000 546.600000 311.200000 ;
      RECT 0.700000 310.400000 546.600000 310.800000 ;
      RECT 0.000000 310.000000 546.600000 310.400000 ;
      RECT 0.700000 309.600000 546.600000 310.000000 ;
      RECT 0.000000 309.200000 546.600000 309.600000 ;
      RECT 0.700000 308.800000 546.600000 309.200000 ;
      RECT 0.000000 308.400000 546.600000 308.800000 ;
      RECT 0.700000 308.000000 546.600000 308.400000 ;
      RECT 0.000000 307.600000 546.600000 308.000000 ;
      RECT 0.700000 307.200000 546.600000 307.600000 ;
      RECT 0.000000 306.800000 546.600000 307.200000 ;
      RECT 0.700000 306.400000 546.600000 306.800000 ;
      RECT 0.000000 306.000000 546.600000 306.400000 ;
      RECT 0.700000 305.600000 546.600000 306.000000 ;
      RECT 0.000000 305.200000 546.600000 305.600000 ;
      RECT 0.700000 304.800000 546.600000 305.200000 ;
      RECT 0.000000 304.400000 546.600000 304.800000 ;
      RECT 0.700000 304.000000 546.600000 304.400000 ;
      RECT 0.000000 303.600000 546.600000 304.000000 ;
      RECT 0.700000 303.200000 546.600000 303.600000 ;
      RECT 0.000000 302.800000 546.600000 303.200000 ;
      RECT 0.700000 302.400000 546.600000 302.800000 ;
      RECT 0.000000 302.000000 546.600000 302.400000 ;
      RECT 0.700000 301.600000 546.600000 302.000000 ;
      RECT 0.000000 301.200000 546.600000 301.600000 ;
      RECT 0.700000 300.800000 546.600000 301.200000 ;
      RECT 0.000000 300.400000 546.600000 300.800000 ;
      RECT 0.700000 300.000000 546.600000 300.400000 ;
      RECT 0.000000 299.600000 546.600000 300.000000 ;
      RECT 0.700000 299.200000 546.600000 299.600000 ;
      RECT 0.000000 298.800000 546.600000 299.200000 ;
      RECT 0.700000 298.400000 546.600000 298.800000 ;
      RECT 0.000000 298.000000 546.600000 298.400000 ;
      RECT 0.700000 297.600000 546.600000 298.000000 ;
      RECT 0.000000 297.200000 546.600000 297.600000 ;
      RECT 0.700000 296.800000 546.600000 297.200000 ;
      RECT 0.000000 296.400000 546.600000 296.800000 ;
      RECT 0.700000 296.000000 546.600000 296.400000 ;
      RECT 0.000000 295.600000 546.600000 296.000000 ;
      RECT 0.700000 295.200000 546.600000 295.600000 ;
      RECT 0.000000 294.800000 546.600000 295.200000 ;
      RECT 0.700000 294.400000 546.600000 294.800000 ;
      RECT 0.000000 294.000000 546.600000 294.400000 ;
      RECT 0.700000 293.600000 546.600000 294.000000 ;
      RECT 0.000000 293.200000 546.600000 293.600000 ;
      RECT 0.700000 292.800000 546.600000 293.200000 ;
      RECT 0.000000 292.400000 546.600000 292.800000 ;
      RECT 0.700000 292.000000 546.600000 292.400000 ;
      RECT 0.000000 291.600000 546.600000 292.000000 ;
      RECT 0.700000 291.200000 546.600000 291.600000 ;
      RECT 0.000000 290.800000 546.600000 291.200000 ;
      RECT 0.700000 290.400000 546.600000 290.800000 ;
      RECT 0.000000 290.000000 546.600000 290.400000 ;
      RECT 0.700000 289.600000 546.600000 290.000000 ;
      RECT 0.000000 289.200000 546.600000 289.600000 ;
      RECT 0.700000 288.800000 546.600000 289.200000 ;
      RECT 0.000000 288.400000 546.600000 288.800000 ;
      RECT 0.700000 288.000000 546.600000 288.400000 ;
      RECT 0.000000 287.600000 546.600000 288.000000 ;
      RECT 0.700000 287.200000 546.600000 287.600000 ;
      RECT 0.000000 286.800000 546.600000 287.200000 ;
      RECT 0.700000 286.400000 546.600000 286.800000 ;
      RECT 0.000000 286.000000 546.600000 286.400000 ;
      RECT 0.700000 285.600000 546.600000 286.000000 ;
      RECT 0.000000 285.200000 546.600000 285.600000 ;
      RECT 0.700000 284.800000 546.600000 285.200000 ;
      RECT 0.000000 284.400000 546.600000 284.800000 ;
      RECT 0.700000 284.000000 546.600000 284.400000 ;
      RECT 0.000000 283.600000 546.600000 284.000000 ;
      RECT 0.700000 283.200000 546.600000 283.600000 ;
      RECT 0.000000 282.800000 546.600000 283.200000 ;
      RECT 0.700000 282.400000 546.600000 282.800000 ;
      RECT 0.000000 282.000000 546.600000 282.400000 ;
      RECT 0.700000 281.600000 546.600000 282.000000 ;
      RECT 0.000000 281.200000 546.600000 281.600000 ;
      RECT 0.700000 280.800000 546.600000 281.200000 ;
      RECT 0.000000 280.400000 546.600000 280.800000 ;
      RECT 0.700000 280.000000 546.600000 280.400000 ;
      RECT 0.000000 279.600000 546.600000 280.000000 ;
      RECT 0.700000 279.200000 546.600000 279.600000 ;
      RECT 0.000000 278.800000 546.600000 279.200000 ;
      RECT 0.700000 278.400000 546.600000 278.800000 ;
      RECT 0.000000 278.000000 546.600000 278.400000 ;
      RECT 0.700000 277.600000 546.600000 278.000000 ;
      RECT 0.000000 277.200000 546.600000 277.600000 ;
      RECT 0.700000 276.800000 546.600000 277.200000 ;
      RECT 0.000000 276.400000 546.600000 276.800000 ;
      RECT 0.700000 276.000000 546.600000 276.400000 ;
      RECT 0.000000 275.600000 546.600000 276.000000 ;
      RECT 0.700000 275.200000 546.600000 275.600000 ;
      RECT 0.000000 274.800000 546.600000 275.200000 ;
      RECT 0.700000 274.400000 546.600000 274.800000 ;
      RECT 0.000000 274.000000 546.600000 274.400000 ;
      RECT 0.700000 273.600000 546.600000 274.000000 ;
      RECT 0.000000 273.200000 546.600000 273.600000 ;
      RECT 0.700000 272.800000 546.600000 273.200000 ;
      RECT 0.000000 272.400000 546.600000 272.800000 ;
      RECT 0.700000 272.000000 546.600000 272.400000 ;
      RECT 0.000000 271.600000 546.600000 272.000000 ;
      RECT 0.700000 271.200000 546.600000 271.600000 ;
      RECT 0.000000 270.800000 546.600000 271.200000 ;
      RECT 0.700000 270.400000 546.600000 270.800000 ;
      RECT 0.000000 270.000000 546.600000 270.400000 ;
      RECT 0.700000 269.600000 546.600000 270.000000 ;
      RECT 0.000000 269.200000 546.600000 269.600000 ;
      RECT 0.700000 268.800000 546.600000 269.200000 ;
      RECT 0.000000 268.400000 546.600000 268.800000 ;
      RECT 0.700000 268.000000 546.600000 268.400000 ;
      RECT 0.000000 267.600000 546.600000 268.000000 ;
      RECT 0.700000 267.200000 546.600000 267.600000 ;
      RECT 0.000000 266.800000 546.600000 267.200000 ;
      RECT 0.700000 266.400000 546.600000 266.800000 ;
      RECT 0.000000 266.000000 546.600000 266.400000 ;
      RECT 0.700000 265.600000 546.600000 266.000000 ;
      RECT 0.000000 265.200000 546.600000 265.600000 ;
      RECT 0.700000 264.800000 546.600000 265.200000 ;
      RECT 0.000000 264.400000 546.600000 264.800000 ;
      RECT 0.700000 264.000000 546.600000 264.400000 ;
      RECT 0.000000 263.600000 546.600000 264.000000 ;
      RECT 0.700000 263.200000 546.600000 263.600000 ;
      RECT 0.000000 262.800000 546.600000 263.200000 ;
      RECT 0.700000 262.400000 546.600000 262.800000 ;
      RECT 0.000000 262.000000 546.600000 262.400000 ;
      RECT 0.700000 261.600000 546.600000 262.000000 ;
      RECT 0.000000 261.200000 546.600000 261.600000 ;
      RECT 0.700000 260.800000 546.600000 261.200000 ;
      RECT 0.000000 260.400000 546.600000 260.800000 ;
      RECT 0.700000 260.000000 546.600000 260.400000 ;
      RECT 0.000000 259.600000 546.600000 260.000000 ;
      RECT 0.700000 259.200000 546.600000 259.600000 ;
      RECT 0.000000 258.800000 546.600000 259.200000 ;
      RECT 0.700000 258.400000 546.600000 258.800000 ;
      RECT 0.000000 258.000000 546.600000 258.400000 ;
      RECT 0.700000 257.600000 546.600000 258.000000 ;
      RECT 0.000000 257.200000 546.600000 257.600000 ;
      RECT 0.700000 256.800000 546.600000 257.200000 ;
      RECT 0.000000 256.400000 546.600000 256.800000 ;
      RECT 0.700000 256.000000 546.600000 256.400000 ;
      RECT 0.000000 255.600000 546.600000 256.000000 ;
      RECT 0.700000 255.200000 546.600000 255.600000 ;
      RECT 0.000000 254.800000 546.600000 255.200000 ;
      RECT 0.700000 254.400000 546.600000 254.800000 ;
      RECT 0.000000 254.000000 546.600000 254.400000 ;
      RECT 0.700000 253.600000 546.600000 254.000000 ;
      RECT 0.000000 253.200000 546.600000 253.600000 ;
      RECT 0.700000 252.800000 546.600000 253.200000 ;
      RECT 0.000000 252.400000 546.600000 252.800000 ;
      RECT 0.700000 252.000000 546.600000 252.400000 ;
      RECT 0.000000 251.600000 546.600000 252.000000 ;
      RECT 0.700000 251.200000 546.600000 251.600000 ;
      RECT 0.000000 250.800000 546.600000 251.200000 ;
      RECT 0.700000 250.400000 546.600000 250.800000 ;
      RECT 0.000000 250.000000 546.600000 250.400000 ;
      RECT 0.700000 249.600000 546.600000 250.000000 ;
      RECT 0.000000 249.200000 546.600000 249.600000 ;
      RECT 0.700000 248.800000 546.600000 249.200000 ;
      RECT 0.000000 248.400000 546.600000 248.800000 ;
      RECT 0.700000 248.000000 546.600000 248.400000 ;
      RECT 0.000000 247.600000 546.600000 248.000000 ;
      RECT 0.700000 247.200000 546.600000 247.600000 ;
      RECT 0.000000 246.800000 546.600000 247.200000 ;
      RECT 0.700000 246.400000 546.600000 246.800000 ;
      RECT 0.000000 246.000000 546.600000 246.400000 ;
      RECT 0.700000 245.600000 546.600000 246.000000 ;
      RECT 0.000000 245.200000 546.600000 245.600000 ;
      RECT 0.700000 244.800000 546.600000 245.200000 ;
      RECT 0.000000 244.400000 546.600000 244.800000 ;
      RECT 0.700000 244.000000 546.600000 244.400000 ;
      RECT 0.000000 243.600000 546.600000 244.000000 ;
      RECT 0.700000 243.200000 546.600000 243.600000 ;
      RECT 0.000000 242.800000 546.600000 243.200000 ;
      RECT 0.700000 242.400000 546.600000 242.800000 ;
      RECT 0.000000 242.000000 546.600000 242.400000 ;
      RECT 0.700000 241.600000 546.600000 242.000000 ;
      RECT 0.000000 241.200000 546.600000 241.600000 ;
      RECT 0.700000 240.800000 546.600000 241.200000 ;
      RECT 0.000000 240.400000 546.600000 240.800000 ;
      RECT 0.700000 240.000000 546.600000 240.400000 ;
      RECT 0.000000 239.600000 546.600000 240.000000 ;
      RECT 0.700000 239.200000 546.600000 239.600000 ;
      RECT 0.000000 238.800000 546.600000 239.200000 ;
      RECT 0.700000 238.400000 546.600000 238.800000 ;
      RECT 0.000000 238.000000 546.600000 238.400000 ;
      RECT 0.700000 237.600000 546.600000 238.000000 ;
      RECT 0.000000 237.200000 546.600000 237.600000 ;
      RECT 0.700000 236.800000 546.600000 237.200000 ;
      RECT 0.000000 236.400000 546.600000 236.800000 ;
      RECT 0.700000 236.000000 546.600000 236.400000 ;
      RECT 0.000000 235.600000 546.600000 236.000000 ;
      RECT 0.700000 235.200000 546.600000 235.600000 ;
      RECT 0.000000 234.800000 546.600000 235.200000 ;
      RECT 0.700000 234.400000 546.600000 234.800000 ;
      RECT 0.000000 234.000000 546.600000 234.400000 ;
      RECT 0.700000 233.600000 546.600000 234.000000 ;
      RECT 0.000000 233.200000 546.600000 233.600000 ;
      RECT 0.700000 232.800000 546.600000 233.200000 ;
      RECT 0.000000 232.400000 546.600000 232.800000 ;
      RECT 0.700000 232.000000 546.600000 232.400000 ;
      RECT 0.000000 231.600000 546.600000 232.000000 ;
      RECT 0.700000 231.200000 546.600000 231.600000 ;
      RECT 0.000000 0.000000 546.600000 231.200000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 546.600000 545.600000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 546.600000 545.600000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 546.600000 545.600000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 546.600000 545.600000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 546.600000 545.600000 ;
  END
END dualcore

END LIBRARY
