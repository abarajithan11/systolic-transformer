##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Wed Mar 22 05:48:36 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO dualcore
  CLASS BLOCK ;
  SIZE 584.600000 BY 583.400000 ;
  FOREIGN dualcore 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 0.150000 0.600000 0.250000 ;
    END
  END clk1
  PIN rst1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 566.150000 0.600000 566.250000 ;
    END
  END rst1
  PIN mem_in_core1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 381.150000 0.600000 381.250000 ;
    END
  END mem_in_core1[31]
  PIN mem_in_core1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 375.550000 0.600000 375.650000 ;
    END
  END mem_in_core1[30]
  PIN mem_in_core1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 369.950000 0.600000 370.050000 ;
    END
  END mem_in_core1[29]
  PIN mem_in_core1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 364.350000 0.600000 364.450000 ;
    END
  END mem_in_core1[28]
  PIN mem_in_core1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 358.750000 0.600000 358.850000 ;
    END
  END mem_in_core1[27]
  PIN mem_in_core1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 353.150000 0.600000 353.250000 ;
    END
  END mem_in_core1[26]
  PIN mem_in_core1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 347.550000 0.600000 347.650000 ;
    END
  END mem_in_core1[25]
  PIN mem_in_core1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 341.950000 0.600000 342.050000 ;
    END
  END mem_in_core1[24]
  PIN mem_in_core1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 336.350000 0.600000 336.450000 ;
    END
  END mem_in_core1[23]
  PIN mem_in_core1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 330.750000 0.600000 330.850000 ;
    END
  END mem_in_core1[22]
  PIN mem_in_core1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 325.150000 0.600000 325.250000 ;
    END
  END mem_in_core1[21]
  PIN mem_in_core1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 319.550000 0.600000 319.650000 ;
    END
  END mem_in_core1[20]
  PIN mem_in_core1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 313.950000 0.600000 314.050000 ;
    END
  END mem_in_core1[19]
  PIN mem_in_core1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 308.350000 0.600000 308.450000 ;
    END
  END mem_in_core1[18]
  PIN mem_in_core1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 302.750000 0.600000 302.850000 ;
    END
  END mem_in_core1[17]
  PIN mem_in_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 297.150000 0.600000 297.250000 ;
    END
  END mem_in_core1[16]
  PIN mem_in_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 291.550000 0.600000 291.650000 ;
    END
  END mem_in_core1[15]
  PIN mem_in_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 285.950000 0.600000 286.050000 ;
    END
  END mem_in_core1[14]
  PIN mem_in_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 280.350000 0.600000 280.450000 ;
    END
  END mem_in_core1[13]
  PIN mem_in_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 274.750000 0.600000 274.850000 ;
    END
  END mem_in_core1[12]
  PIN mem_in_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 269.150000 0.600000 269.250000 ;
    END
  END mem_in_core1[11]
  PIN mem_in_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 263.550000 0.600000 263.650000 ;
    END
  END mem_in_core1[10]
  PIN mem_in_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 257.950000 0.600000 258.050000 ;
    END
  END mem_in_core1[9]
  PIN mem_in_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 252.350000 0.600000 252.450000 ;
    END
  END mem_in_core1[8]
  PIN mem_in_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 246.750000 0.600000 246.850000 ;
    END
  END mem_in_core1[7]
  PIN mem_in_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 241.150000 0.600000 241.250000 ;
    END
  END mem_in_core1[6]
  PIN mem_in_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 235.550000 0.600000 235.650000 ;
    END
  END mem_in_core1[5]
  PIN mem_in_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 229.950000 0.600000 230.050000 ;
    END
  END mem_in_core1[4]
  PIN mem_in_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 224.350000 0.600000 224.450000 ;
    END
  END mem_in_core1[3]
  PIN mem_in_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 218.750000 0.600000 218.850000 ;
    END
  END mem_in_core1[2]
  PIN mem_in_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 213.150000 0.600000 213.250000 ;
    END
  END mem_in_core1[1]
  PIN mem_in_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 207.550000 0.600000 207.650000 ;
    END
  END mem_in_core1[0]
  PIN inst_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 106.550000 0.600000 106.650000 ;
    END
  END inst_core1[16]
  PIN inst_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 100.950000 0.600000 101.050000 ;
    END
  END inst_core1[15]
  PIN inst_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 95.350000 0.600000 95.450000 ;
    END
  END inst_core1[14]
  PIN inst_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 89.750000 0.600000 89.850000 ;
    END
  END inst_core1[13]
  PIN inst_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 84.150000 0.600000 84.250000 ;
    END
  END inst_core1[12]
  PIN inst_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 78.550000 0.600000 78.650000 ;
    END
  END inst_core1[11]
  PIN inst_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 72.950000 0.600000 73.050000 ;
    END
  END inst_core1[10]
  PIN inst_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 67.350000 0.600000 67.450000 ;
    END
  END inst_core1[9]
  PIN inst_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 61.750000 0.600000 61.850000 ;
    END
  END inst_core1[8]
  PIN inst_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 56.150000 0.600000 56.250000 ;
    END
  END inst_core1[7]
  PIN inst_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 50.550000 0.600000 50.650000 ;
    END
  END inst_core1[6]
  PIN inst_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 44.950000 0.600000 45.050000 ;
    END
  END inst_core1[5]
  PIN inst_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 39.350000 0.600000 39.450000 ;
    END
  END inst_core1[4]
  PIN inst_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 33.750000 0.600000 33.850000 ;
    END
  END inst_core1[3]
  PIN inst_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 28.150000 0.600000 28.250000 ;
    END
  END inst_core1[2]
  PIN inst_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 22.550000 0.600000 22.650000 ;
    END
  END inst_core1[1]
  PIN inst_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 16.950000 0.600000 17.050000 ;
    END
  END inst_core1[0]
  PIN out_core1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 259.650000 0.000000 259.750000 0.600000 ;
    END
  END out_core1[87]
  PIN out_core1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 256.650000 0.000000 256.750000 0.600000 ;
    END
  END out_core1[86]
  PIN out_core1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 253.850000 0.000000 253.950000 0.600000 ;
    END
  END out_core1[85]
  PIN out_core1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 250.850000 0.000000 250.950000 0.600000 ;
    END
  END out_core1[84]
  PIN out_core1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 247.850000 0.000000 247.950000 0.600000 ;
    END
  END out_core1[83]
  PIN out_core1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 244.850000 0.000000 244.950000 0.600000 ;
    END
  END out_core1[82]
  PIN out_core1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 242.050000 0.000000 242.150000 0.600000 ;
    END
  END out_core1[81]
  PIN out_core1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 239.050000 0.000000 239.150000 0.600000 ;
    END
  END out_core1[80]
  PIN out_core1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 236.050000 0.000000 236.150000 0.600000 ;
    END
  END out_core1[79]
  PIN out_core1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 233.050000 0.000000 233.150000 0.600000 ;
    END
  END out_core1[78]
  PIN out_core1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 230.250000 0.000000 230.350000 0.600000 ;
    END
  END out_core1[77]
  PIN out_core1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 227.250000 0.000000 227.350000 0.600000 ;
    END
  END out_core1[76]
  PIN out_core1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 224.250000 0.000000 224.350000 0.600000 ;
    END
  END out_core1[75]
  PIN out_core1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.250000 0.000000 221.350000 0.600000 ;
    END
  END out_core1[74]
  PIN out_core1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 218.450000 0.000000 218.550000 0.600000 ;
    END
  END out_core1[73]
  PIN out_core1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.450000 0.000000 215.550000 0.600000 ;
    END
  END out_core1[72]
  PIN out_core1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 212.450000 0.000000 212.550000 0.600000 ;
    END
  END out_core1[71]
  PIN out_core1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.450000 0.000000 209.550000 0.600000 ;
    END
  END out_core1[70]
  PIN out_core1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 206.650000 0.000000 206.750000 0.600000 ;
    END
  END out_core1[69]
  PIN out_core1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 203.650000 0.000000 203.750000 0.600000 ;
    END
  END out_core1[68]
  PIN out_core1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 200.650000 0.000000 200.750000 0.600000 ;
    END
  END out_core1[67]
  PIN out_core1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.650000 0.000000 197.750000 0.600000 ;
    END
  END out_core1[66]
  PIN out_core1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 194.650000 0.000000 194.750000 0.600000 ;
    END
  END out_core1[65]
  PIN out_core1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.850000 0.000000 191.950000 0.600000 ;
    END
  END out_core1[64]
  PIN out_core1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 188.850000 0.000000 188.950000 0.600000 ;
    END
  END out_core1[63]
  PIN out_core1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.850000 0.000000 185.950000 0.600000 ;
    END
  END out_core1[62]
  PIN out_core1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 182.850000 0.000000 182.950000 0.600000 ;
    END
  END out_core1[61]
  PIN out_core1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.050000 0.000000 180.150000 0.600000 ;
    END
  END out_core1[60]
  PIN out_core1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.050000 0.000000 177.150000 0.600000 ;
    END
  END out_core1[59]
  PIN out_core1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 174.050000 0.000000 174.150000 0.600000 ;
    END
  END out_core1[58]
  PIN out_core1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 171.050000 0.000000 171.150000 0.600000 ;
    END
  END out_core1[57]
  PIN out_core1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.250000 0.000000 168.350000 0.600000 ;
    END
  END out_core1[56]
  PIN out_core1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.250000 0.000000 165.350000 0.600000 ;
    END
  END out_core1[55]
  PIN out_core1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.250000 0.000000 162.350000 0.600000 ;
    END
  END out_core1[54]
  PIN out_core1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.250000 0.000000 159.350000 0.600000 ;
    END
  END out_core1[53]
  PIN out_core1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.450000 0.000000 156.550000 0.600000 ;
    END
  END out_core1[52]
  PIN out_core1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.450000 0.000000 153.550000 0.600000 ;
    END
  END out_core1[51]
  PIN out_core1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 150.450000 0.000000 150.550000 0.600000 ;
    END
  END out_core1[50]
  PIN out_core1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 147.450000 0.000000 147.550000 0.600000 ;
    END
  END out_core1[49]
  PIN out_core1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 144.650000 0.000000 144.750000 0.600000 ;
    END
  END out_core1[48]
  PIN out_core1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.650000 0.000000 141.750000 0.600000 ;
    END
  END out_core1[47]
  PIN out_core1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.650000 0.000000 138.750000 0.600000 ;
    END
  END out_core1[46]
  PIN out_core1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.650000 0.000000 135.750000 0.600000 ;
    END
  END out_core1[45]
  PIN out_core1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.850000 0.000000 132.950000 0.600000 ;
    END
  END out_core1[44]
  PIN out_core1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.850000 0.000000 129.950000 0.600000 ;
    END
  END out_core1[43]
  PIN out_core1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 126.850000 0.000000 126.950000 0.600000 ;
    END
  END out_core1[42]
  PIN out_core1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 123.850000 0.000000 123.950000 0.600000 ;
    END
  END out_core1[41]
  PIN out_core1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.050000 0.000000 121.150000 0.600000 ;
    END
  END out_core1[40]
  PIN out_core1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 118.050000 0.000000 118.150000 0.600000 ;
    END
  END out_core1[39]
  PIN out_core1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 115.050000 0.000000 115.150000 0.600000 ;
    END
  END out_core1[38]
  PIN out_core1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 112.050000 0.000000 112.150000 0.600000 ;
    END
  END out_core1[37]
  PIN out_core1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.250000 0.000000 109.350000 0.600000 ;
    END
  END out_core1[36]
  PIN out_core1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.250000 0.000000 106.350000 0.600000 ;
    END
  END out_core1[35]
  PIN out_core1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.250000 0.000000 103.350000 0.600000 ;
    END
  END out_core1[34]
  PIN out_core1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.250000 0.000000 100.350000 0.600000 ;
    END
  END out_core1[33]
  PIN out_core1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.250000 0.000000 97.350000 0.600000 ;
    END
  END out_core1[32]
  PIN out_core1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 94.450000 0.000000 94.550000 0.600000 ;
    END
  END out_core1[31]
  PIN out_core1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 91.450000 0.000000 91.550000 0.600000 ;
    END
  END out_core1[30]
  PIN out_core1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 88.450000 0.000000 88.550000 0.600000 ;
    END
  END out_core1[29]
  PIN out_core1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.450000 0.000000 85.550000 0.600000 ;
    END
  END out_core1[28]
  PIN out_core1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.650000 0.000000 82.750000 0.600000 ;
    END
  END out_core1[27]
  PIN out_core1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.650000 0.000000 79.750000 0.600000 ;
    END
  END out_core1[26]
  PIN out_core1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.650000 0.000000 76.750000 0.600000 ;
    END
  END out_core1[25]
  PIN out_core1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.650000 0.000000 73.750000 0.600000 ;
    END
  END out_core1[24]
  PIN out_core1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 70.850000 0.000000 70.950000 0.600000 ;
    END
  END out_core1[23]
  PIN out_core1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 67.850000 0.000000 67.950000 0.600000 ;
    END
  END out_core1[22]
  PIN out_core1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 64.850000 0.000000 64.950000 0.600000 ;
    END
  END out_core1[21]
  PIN out_core1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 61.850000 0.000000 61.950000 0.600000 ;
    END
  END out_core1[20]
  PIN out_core1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 59.050000 0.000000 59.150000 0.600000 ;
    END
  END out_core1[19]
  PIN out_core1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 56.050000 0.000000 56.150000 0.600000 ;
    END
  END out_core1[18]
  PIN out_core1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 53.050000 0.000000 53.150000 0.600000 ;
    END
  END out_core1[17]
  PIN out_core1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 50.050000 0.000000 50.150000 0.600000 ;
    END
  END out_core1[16]
  PIN out_core1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 47.250000 0.000000 47.350000 0.600000 ;
    END
  END out_core1[15]
  PIN out_core1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 44.250000 0.000000 44.350000 0.600000 ;
    END
  END out_core1[14]
  PIN out_core1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 41.250000 0.000000 41.350000 0.600000 ;
    END
  END out_core1[13]
  PIN out_core1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 38.250000 0.000000 38.350000 0.600000 ;
    END
  END out_core1[12]
  PIN out_core1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 35.450000 0.000000 35.550000 0.600000 ;
    END
  END out_core1[11]
  PIN out_core1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 32.450000 0.000000 32.550000 0.600000 ;
    END
  END out_core1[10]
  PIN out_core1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 29.450000 0.000000 29.550000 0.600000 ;
    END
  END out_core1[9]
  PIN out_core1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 26.450000 0.000000 26.550000 0.600000 ;
    END
  END out_core1[8]
  PIN out_core1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 23.650000 0.000000 23.750000 0.600000 ;
    END
  END out_core1[7]
  PIN out_core1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 20.650000 0.000000 20.750000 0.600000 ;
    END
  END out_core1[6]
  PIN out_core1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 17.650000 0.000000 17.750000 0.600000 ;
    END
  END out_core1[5]
  PIN out_core1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 14.650000 0.000000 14.750000 0.600000 ;
    END
  END out_core1[4]
  PIN out_core1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 11.850000 0.000000 11.950000 0.600000 ;
    END
  END out_core1[3]
  PIN out_core1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 8.850000 0.000000 8.950000 0.600000 ;
    END
  END out_core1[2]
  PIN out_core1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5.850000 0.000000 5.950000 0.600000 ;
    END
  END out_core1[1]
  PIN out_core1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.850000 0.000000 2.950000 0.600000 ;
    END
  END out_core1[0]
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 5.750000 0.600000 5.850000 ;
    END
  END clk2
  PIN rst2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 571.750000 0.600000 571.850000 ;
    END
  END rst2
  PIN mem_in_core2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 560.550000 0.600000 560.650000 ;
    END
  END mem_in_core2[31]
  PIN mem_in_core2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 554.950000 0.600000 555.050000 ;
    END
  END mem_in_core2[30]
  PIN mem_in_core2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 549.350000 0.600000 549.450000 ;
    END
  END mem_in_core2[29]
  PIN mem_in_core2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 543.750000 0.600000 543.850000 ;
    END
  END mem_in_core2[28]
  PIN mem_in_core2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 538.150000 0.600000 538.250000 ;
    END
  END mem_in_core2[27]
  PIN mem_in_core2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 532.550000 0.600000 532.650000 ;
    END
  END mem_in_core2[26]
  PIN mem_in_core2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 526.950000 0.600000 527.050000 ;
    END
  END mem_in_core2[25]
  PIN mem_in_core2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 521.350000 0.600000 521.450000 ;
    END
  END mem_in_core2[24]
  PIN mem_in_core2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 515.750000 0.600000 515.850000 ;
    END
  END mem_in_core2[23]
  PIN mem_in_core2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 510.150000 0.600000 510.250000 ;
    END
  END mem_in_core2[22]
  PIN mem_in_core2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 504.550000 0.600000 504.650000 ;
    END
  END mem_in_core2[21]
  PIN mem_in_core2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 498.950000 0.600000 499.050000 ;
    END
  END mem_in_core2[20]
  PIN mem_in_core2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 493.350000 0.600000 493.450000 ;
    END
  END mem_in_core2[19]
  PIN mem_in_core2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 487.750000 0.600000 487.850000 ;
    END
  END mem_in_core2[18]
  PIN mem_in_core2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 482.150000 0.600000 482.250000 ;
    END
  END mem_in_core2[17]
  PIN mem_in_core2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 476.550000 0.600000 476.650000 ;
    END
  END mem_in_core2[16]
  PIN mem_in_core2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 470.950000 0.600000 471.050000 ;
    END
  END mem_in_core2[15]
  PIN mem_in_core2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 465.350000 0.600000 465.450000 ;
    END
  END mem_in_core2[14]
  PIN mem_in_core2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 459.750000 0.600000 459.850000 ;
    END
  END mem_in_core2[13]
  PIN mem_in_core2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 454.150000 0.600000 454.250000 ;
    END
  END mem_in_core2[12]
  PIN mem_in_core2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 448.550000 0.600000 448.650000 ;
    END
  END mem_in_core2[11]
  PIN mem_in_core2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 442.950000 0.600000 443.050000 ;
    END
  END mem_in_core2[10]
  PIN mem_in_core2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 437.350000 0.600000 437.450000 ;
    END
  END mem_in_core2[9]
  PIN mem_in_core2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 431.750000 0.600000 431.850000 ;
    END
  END mem_in_core2[8]
  PIN mem_in_core2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 426.150000 0.600000 426.250000 ;
    END
  END mem_in_core2[7]
  PIN mem_in_core2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 420.550000 0.600000 420.650000 ;
    END
  END mem_in_core2[6]
  PIN mem_in_core2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 414.950000 0.600000 415.050000 ;
    END
  END mem_in_core2[5]
  PIN mem_in_core2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 409.350000 0.600000 409.450000 ;
    END
  END mem_in_core2[4]
  PIN mem_in_core2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 403.750000 0.600000 403.850000 ;
    END
  END mem_in_core2[3]
  PIN mem_in_core2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 398.150000 0.600000 398.250000 ;
    END
  END mem_in_core2[2]
  PIN mem_in_core2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 392.550000 0.600000 392.650000 ;
    END
  END mem_in_core2[1]
  PIN mem_in_core2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 386.750000 0.600000 386.850000 ;
    END
  END mem_in_core2[0]
  PIN inst_core2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 201.950000 0.600000 202.050000 ;
    END
  END inst_core2[16]
  PIN inst_core2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 196.350000 0.600000 196.450000 ;
    END
  END inst_core2[15]
  PIN inst_core2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 190.550000 0.600000 190.650000 ;
    END
  END inst_core2[14]
  PIN inst_core2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 184.950000 0.600000 185.050000 ;
    END
  END inst_core2[13]
  PIN inst_core2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 179.350000 0.600000 179.450000 ;
    END
  END inst_core2[12]
  PIN inst_core2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 173.750000 0.600000 173.850000 ;
    END
  END inst_core2[11]
  PIN inst_core2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 168.150000 0.600000 168.250000 ;
    END
  END inst_core2[10]
  PIN inst_core2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 162.550000 0.600000 162.650000 ;
    END
  END inst_core2[9]
  PIN inst_core2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 156.950000 0.600000 157.050000 ;
    END
  END inst_core2[8]
  PIN inst_core2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 151.350000 0.600000 151.450000 ;
    END
  END inst_core2[7]
  PIN inst_core2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 145.750000 0.600000 145.850000 ;
    END
  END inst_core2[6]
  PIN inst_core2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 140.150000 0.600000 140.250000 ;
    END
  END inst_core2[5]
  PIN inst_core2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 134.550000 0.600000 134.650000 ;
    END
  END inst_core2[4]
  PIN inst_core2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 128.950000 0.600000 129.050000 ;
    END
  END inst_core2[3]
  PIN inst_core2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 123.350000 0.600000 123.450000 ;
    END
  END inst_core2[2]
  PIN inst_core2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 117.750000 0.600000 117.850000 ;
    END
  END inst_core2[1]
  PIN inst_core2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 112.150000 0.600000 112.250000 ;
    END
  END inst_core2[0]
  PIN out_core2[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 519.450000 0.000000 519.550000 0.600000 ;
    END
  END out_core2[87]
  PIN out_core2[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 516.450000 0.000000 516.550000 0.600000 ;
    END
  END out_core2[86]
  PIN out_core2[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 513.450000 0.000000 513.550000 0.600000 ;
    END
  END out_core2[85]
  PIN out_core2[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 510.650000 0.000000 510.750000 0.600000 ;
    END
  END out_core2[84]
  PIN out_core2[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 507.650000 0.000000 507.750000 0.600000 ;
    END
  END out_core2[83]
  PIN out_core2[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 504.650000 0.000000 504.750000 0.600000 ;
    END
  END out_core2[82]
  PIN out_core2[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 501.650000 0.000000 501.750000 0.600000 ;
    END
  END out_core2[81]
  PIN out_core2[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 498.850000 0.000000 498.950000 0.600000 ;
    END
  END out_core2[80]
  PIN out_core2[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 495.850000 0.000000 495.950000 0.600000 ;
    END
  END out_core2[79]
  PIN out_core2[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 492.850000 0.000000 492.950000 0.600000 ;
    END
  END out_core2[78]
  PIN out_core2[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 489.850000 0.000000 489.950000 0.600000 ;
    END
  END out_core2[77]
  PIN out_core2[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 487.050000 0.000000 487.150000 0.600000 ;
    END
  END out_core2[76]
  PIN out_core2[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 484.050000 0.000000 484.150000 0.600000 ;
    END
  END out_core2[75]
  PIN out_core2[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 481.050000 0.000000 481.150000 0.600000 ;
    END
  END out_core2[74]
  PIN out_core2[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 478.050000 0.000000 478.150000 0.600000 ;
    END
  END out_core2[73]
  PIN out_core2[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 475.050000 0.000000 475.150000 0.600000 ;
    END
  END out_core2[72]
  PIN out_core2[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 472.250000 0.000000 472.350000 0.600000 ;
    END
  END out_core2[71]
  PIN out_core2[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 469.250000 0.000000 469.350000 0.600000 ;
    END
  END out_core2[70]
  PIN out_core2[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 466.250000 0.000000 466.350000 0.600000 ;
    END
  END out_core2[69]
  PIN out_core2[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 463.250000 0.000000 463.350000 0.600000 ;
    END
  END out_core2[68]
  PIN out_core2[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 460.450000 0.000000 460.550000 0.600000 ;
    END
  END out_core2[67]
  PIN out_core2[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 457.450000 0.000000 457.550000 0.600000 ;
    END
  END out_core2[66]
  PIN out_core2[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 454.450000 0.000000 454.550000 0.600000 ;
    END
  END out_core2[65]
  PIN out_core2[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 451.450000 0.000000 451.550000 0.600000 ;
    END
  END out_core2[64]
  PIN out_core2[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 448.650000 0.000000 448.750000 0.600000 ;
    END
  END out_core2[63]
  PIN out_core2[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 445.650000 0.000000 445.750000 0.600000 ;
    END
  END out_core2[62]
  PIN out_core2[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 442.650000 0.000000 442.750000 0.600000 ;
    END
  END out_core2[61]
  PIN out_core2[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 439.650000 0.000000 439.750000 0.600000 ;
    END
  END out_core2[60]
  PIN out_core2[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 436.850000 0.000000 436.950000 0.600000 ;
    END
  END out_core2[59]
  PIN out_core2[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 433.850000 0.000000 433.950000 0.600000 ;
    END
  END out_core2[58]
  PIN out_core2[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 430.850000 0.000000 430.950000 0.600000 ;
    END
  END out_core2[57]
  PIN out_core2[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 427.850000 0.000000 427.950000 0.600000 ;
    END
  END out_core2[56]
  PIN out_core2[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 425.050000 0.000000 425.150000 0.600000 ;
    END
  END out_core2[55]
  PIN out_core2[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 422.050000 0.000000 422.150000 0.600000 ;
    END
  END out_core2[54]
  PIN out_core2[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 419.050000 0.000000 419.150000 0.600000 ;
    END
  END out_core2[53]
  PIN out_core2[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 416.050000 0.000000 416.150000 0.600000 ;
    END
  END out_core2[52]
  PIN out_core2[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 413.250000 0.000000 413.350000 0.600000 ;
    END
  END out_core2[51]
  PIN out_core2[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 410.250000 0.000000 410.350000 0.600000 ;
    END
  END out_core2[50]
  PIN out_core2[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 407.250000 0.000000 407.350000 0.600000 ;
    END
  END out_core2[49]
  PIN out_core2[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 404.250000 0.000000 404.350000 0.600000 ;
    END
  END out_core2[48]
  PIN out_core2[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.450000 0.000000 401.550000 0.600000 ;
    END
  END out_core2[47]
  PIN out_core2[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 398.450000 0.000000 398.550000 0.600000 ;
    END
  END out_core2[46]
  PIN out_core2[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 395.450000 0.000000 395.550000 0.600000 ;
    END
  END out_core2[45]
  PIN out_core2[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 392.450000 0.000000 392.550000 0.600000 ;
    END
  END out_core2[44]
  PIN out_core2[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 389.450000 0.000000 389.550000 0.600000 ;
    END
  END out_core2[43]
  PIN out_core2[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 386.650000 0.000000 386.750000 0.600000 ;
    END
  END out_core2[42]
  PIN out_core2[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 383.650000 0.000000 383.750000 0.600000 ;
    END
  END out_core2[41]
  PIN out_core2[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380.650000 0.000000 380.750000 0.600000 ;
    END
  END out_core2[40]
  PIN out_core2[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 377.650000 0.000000 377.750000 0.600000 ;
    END
  END out_core2[39]
  PIN out_core2[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 374.850000 0.000000 374.950000 0.600000 ;
    END
  END out_core2[38]
  PIN out_core2[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 371.850000 0.000000 371.950000 0.600000 ;
    END
  END out_core2[37]
  PIN out_core2[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 368.850000 0.000000 368.950000 0.600000 ;
    END
  END out_core2[36]
  PIN out_core2[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 365.850000 0.000000 365.950000 0.600000 ;
    END
  END out_core2[35]
  PIN out_core2[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 363.050000 0.000000 363.150000 0.600000 ;
    END
  END out_core2[34]
  PIN out_core2[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 360.050000 0.000000 360.150000 0.600000 ;
    END
  END out_core2[33]
  PIN out_core2[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 357.050000 0.000000 357.150000 0.600000 ;
    END
  END out_core2[32]
  PIN out_core2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 354.050000 0.000000 354.150000 0.600000 ;
    END
  END out_core2[31]
  PIN out_core2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 351.250000 0.000000 351.350000 0.600000 ;
    END
  END out_core2[30]
  PIN out_core2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 348.250000 0.000000 348.350000 0.600000 ;
    END
  END out_core2[29]
  PIN out_core2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 345.250000 0.000000 345.350000 0.600000 ;
    END
  END out_core2[28]
  PIN out_core2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 342.250000 0.000000 342.350000 0.600000 ;
    END
  END out_core2[27]
  PIN out_core2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 339.450000 0.000000 339.550000 0.600000 ;
    END
  END out_core2[26]
  PIN out_core2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 336.450000 0.000000 336.550000 0.600000 ;
    END
  END out_core2[25]
  PIN out_core2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 333.450000 0.000000 333.550000 0.600000 ;
    END
  END out_core2[24]
  PIN out_core2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 330.450000 0.000000 330.550000 0.600000 ;
    END
  END out_core2[23]
  PIN out_core2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.650000 0.000000 327.750000 0.600000 ;
    END
  END out_core2[22]
  PIN out_core2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 324.650000 0.000000 324.750000 0.600000 ;
    END
  END out_core2[21]
  PIN out_core2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 321.650000 0.000000 321.750000 0.600000 ;
    END
  END out_core2[20]
  PIN out_core2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 318.650000 0.000000 318.750000 0.600000 ;
    END
  END out_core2[19]
  PIN out_core2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 315.850000 0.000000 315.950000 0.600000 ;
    END
  END out_core2[18]
  PIN out_core2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 312.850000 0.000000 312.950000 0.600000 ;
    END
  END out_core2[17]
  PIN out_core2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 309.850000 0.000000 309.950000 0.600000 ;
    END
  END out_core2[16]
  PIN out_core2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 306.850000 0.000000 306.950000 0.600000 ;
    END
  END out_core2[15]
  PIN out_core2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 304.050000 0.000000 304.150000 0.600000 ;
    END
  END out_core2[14]
  PIN out_core2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 301.050000 0.000000 301.150000 0.600000 ;
    END
  END out_core2[13]
  PIN out_core2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.050000 0.000000 298.150000 0.600000 ;
    END
  END out_core2[12]
  PIN out_core2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.050000 0.000000 295.150000 0.600000 ;
    END
  END out_core2[11]
  PIN out_core2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 292.050000 0.000000 292.150000 0.600000 ;
    END
  END out_core2[10]
  PIN out_core2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 289.250000 0.000000 289.350000 0.600000 ;
    END
  END out_core2[9]
  PIN out_core2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 286.250000 0.000000 286.350000 0.600000 ;
    END
  END out_core2[8]
  PIN out_core2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 283.250000 0.000000 283.350000 0.600000 ;
    END
  END out_core2[7]
  PIN out_core2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 280.250000 0.000000 280.350000 0.600000 ;
    END
  END out_core2[6]
  PIN out_core2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 277.450000 0.000000 277.550000 0.600000 ;
    END
  END out_core2[5]
  PIN out_core2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 274.450000 0.000000 274.550000 0.600000 ;
    END
  END out_core2[4]
  PIN out_core2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 271.450000 0.000000 271.550000 0.600000 ;
    END
  END out_core2[3]
  PIN out_core2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 268.450000 0.000000 268.550000 0.600000 ;
    END
  END out_core2[2]
  PIN out_core2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 265.650000 0.000000 265.750000 0.600000 ;
    END
  END out_core2[1]
  PIN out_core2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 262.650000 0.000000 262.750000 0.600000 ;
    END
  END out_core2[0]
  PIN norm_gate
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 11.350000 0.600000 11.450000 ;
    END
  END norm_gate
  PIN s_valid1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 577.350000 0.600000 577.450000 ;
    END
  END s_valid1
  PIN s_valid2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 583.150000 0.600000 583.250000 ;
    END
  END s_valid2
  PIN psum_norm_1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 551.850000 0.000000 551.950000 0.600000 ;
    END
  END psum_norm_1[10]
  PIN psum_norm_1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 548.850000 0.000000 548.950000 0.600000 ;
    END
  END psum_norm_1[9]
  PIN psum_norm_1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 546.050000 0.000000 546.150000 0.600000 ;
    END
  END psum_norm_1[8]
  PIN psum_norm_1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 543.050000 0.000000 543.150000 0.600000 ;
    END
  END psum_norm_1[7]
  PIN psum_norm_1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 540.050000 0.000000 540.150000 0.600000 ;
    END
  END psum_norm_1[6]
  PIN psum_norm_1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 537.050000 0.000000 537.150000 0.600000 ;
    END
  END psum_norm_1[5]
  PIN psum_norm_1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 534.250000 0.000000 534.350000 0.600000 ;
    END
  END psum_norm_1[4]
  PIN psum_norm_1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 531.250000 0.000000 531.350000 0.600000 ;
    END
  END psum_norm_1[3]
  PIN psum_norm_1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 528.250000 0.000000 528.350000 0.600000 ;
    END
  END psum_norm_1[2]
  PIN psum_norm_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 525.250000 0.000000 525.350000 0.600000 ;
    END
  END psum_norm_1[1]
  PIN psum_norm_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 522.450000 0.000000 522.550000 0.600000 ;
    END
  END psum_norm_1[0]
  PIN psum_norm_2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 584.450000 0.000000 584.550000 0.600000 ;
    END
  END psum_norm_2[10]
  PIN psum_norm_2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 581.450000 0.000000 581.550000 0.600000 ;
    END
  END psum_norm_2[9]
  PIN psum_norm_2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 578.450000 0.000000 578.550000 0.600000 ;
    END
  END psum_norm_2[8]
  PIN psum_norm_2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 575.450000 0.000000 575.550000 0.600000 ;
    END
  END psum_norm_2[7]
  PIN psum_norm_2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 572.450000 0.000000 572.550000 0.600000 ;
    END
  END psum_norm_2[6]
  PIN psum_norm_2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 569.650000 0.000000 569.750000 0.600000 ;
    END
  END psum_norm_2[5]
  PIN psum_norm_2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 566.650000 0.000000 566.750000 0.600000 ;
    END
  END psum_norm_2[4]
  PIN psum_norm_2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 563.650000 0.000000 563.750000 0.600000 ;
    END
  END psum_norm_2[3]
  PIN psum_norm_2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 560.650000 0.000000 560.750000 0.600000 ;
    END
  END psum_norm_2[2]
  PIN psum_norm_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 557.850000 0.000000 557.950000 0.600000 ;
    END
  END psum_norm_2[1]
  PIN psum_norm_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 554.850000 0.000000 554.950000 0.600000 ;
    END
  END psum_norm_2[0]
  PIN norm_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.850000 0.000000 0.950000 0.600000 ;
    END
  END norm_valid
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 584.600000 583.400000 ;
    LAYER M2 ;
      RECT 0.000000 0.000000 584.600000 583.400000 ;
    LAYER M3 ;
      RECT 0.000000 583.350000 584.600000 583.400000 ;
      RECT 0.720000 583.050000 584.600000 583.350000 ;
      RECT 0.000000 577.550000 584.600000 583.050000 ;
      RECT 0.720000 577.250000 584.600000 577.550000 ;
      RECT 0.000000 571.950000 584.600000 577.250000 ;
      RECT 0.720000 571.650000 584.600000 571.950000 ;
      RECT 0.000000 566.350000 584.600000 571.650000 ;
      RECT 0.720000 566.050000 584.600000 566.350000 ;
      RECT 0.000000 560.750000 584.600000 566.050000 ;
      RECT 0.720000 560.450000 584.600000 560.750000 ;
      RECT 0.000000 555.150000 584.600000 560.450000 ;
      RECT 0.720000 554.850000 584.600000 555.150000 ;
      RECT 0.000000 549.550000 584.600000 554.850000 ;
      RECT 0.720000 549.250000 584.600000 549.550000 ;
      RECT 0.000000 543.950000 584.600000 549.250000 ;
      RECT 0.720000 543.650000 584.600000 543.950000 ;
      RECT 0.000000 538.350000 584.600000 543.650000 ;
      RECT 0.720000 538.050000 584.600000 538.350000 ;
      RECT 0.000000 532.750000 584.600000 538.050000 ;
      RECT 0.720000 532.450000 584.600000 532.750000 ;
      RECT 0.000000 527.150000 584.600000 532.450000 ;
      RECT 0.720000 526.850000 584.600000 527.150000 ;
      RECT 0.000000 521.550000 584.600000 526.850000 ;
      RECT 0.720000 521.250000 584.600000 521.550000 ;
      RECT 0.000000 515.950000 584.600000 521.250000 ;
      RECT 0.720000 515.650000 584.600000 515.950000 ;
      RECT 0.000000 510.350000 584.600000 515.650000 ;
      RECT 0.720000 510.050000 584.600000 510.350000 ;
      RECT 0.000000 504.750000 584.600000 510.050000 ;
      RECT 0.720000 504.450000 584.600000 504.750000 ;
      RECT 0.000000 499.150000 584.600000 504.450000 ;
      RECT 0.720000 498.850000 584.600000 499.150000 ;
      RECT 0.000000 493.550000 584.600000 498.850000 ;
      RECT 0.720000 493.250000 584.600000 493.550000 ;
      RECT 0.000000 487.950000 584.600000 493.250000 ;
      RECT 0.720000 487.650000 584.600000 487.950000 ;
      RECT 0.000000 482.350000 584.600000 487.650000 ;
      RECT 0.720000 482.050000 584.600000 482.350000 ;
      RECT 0.000000 476.750000 584.600000 482.050000 ;
      RECT 0.720000 476.450000 584.600000 476.750000 ;
      RECT 0.000000 471.150000 584.600000 476.450000 ;
      RECT 0.720000 470.850000 584.600000 471.150000 ;
      RECT 0.000000 465.550000 584.600000 470.850000 ;
      RECT 0.720000 465.250000 584.600000 465.550000 ;
      RECT 0.000000 459.950000 584.600000 465.250000 ;
      RECT 0.720000 459.650000 584.600000 459.950000 ;
      RECT 0.000000 454.350000 584.600000 459.650000 ;
      RECT 0.720000 454.050000 584.600000 454.350000 ;
      RECT 0.000000 448.750000 584.600000 454.050000 ;
      RECT 0.720000 448.450000 584.600000 448.750000 ;
      RECT 0.000000 443.150000 584.600000 448.450000 ;
      RECT 0.720000 442.850000 584.600000 443.150000 ;
      RECT 0.000000 437.550000 584.600000 442.850000 ;
      RECT 0.720000 437.250000 584.600000 437.550000 ;
      RECT 0.000000 431.950000 584.600000 437.250000 ;
      RECT 0.720000 431.650000 584.600000 431.950000 ;
      RECT 0.000000 426.350000 584.600000 431.650000 ;
      RECT 0.720000 426.050000 584.600000 426.350000 ;
      RECT 0.000000 420.750000 584.600000 426.050000 ;
      RECT 0.720000 420.450000 584.600000 420.750000 ;
      RECT 0.000000 415.150000 584.600000 420.450000 ;
      RECT 0.720000 414.850000 584.600000 415.150000 ;
      RECT 0.000000 409.550000 584.600000 414.850000 ;
      RECT 0.720000 409.250000 584.600000 409.550000 ;
      RECT 0.000000 403.950000 584.600000 409.250000 ;
      RECT 0.720000 403.650000 584.600000 403.950000 ;
      RECT 0.000000 398.350000 584.600000 403.650000 ;
      RECT 0.720000 398.050000 584.600000 398.350000 ;
      RECT 0.000000 392.750000 584.600000 398.050000 ;
      RECT 0.720000 392.450000 584.600000 392.750000 ;
      RECT 0.000000 386.950000 584.600000 392.450000 ;
      RECT 0.720000 386.650000 584.600000 386.950000 ;
      RECT 0.000000 381.350000 584.600000 386.650000 ;
      RECT 0.720000 381.050000 584.600000 381.350000 ;
      RECT 0.000000 375.750000 584.600000 381.050000 ;
      RECT 0.720000 375.450000 584.600000 375.750000 ;
      RECT 0.000000 370.150000 584.600000 375.450000 ;
      RECT 0.720000 369.850000 584.600000 370.150000 ;
      RECT 0.000000 364.550000 584.600000 369.850000 ;
      RECT 0.720000 364.250000 584.600000 364.550000 ;
      RECT 0.000000 358.950000 584.600000 364.250000 ;
      RECT 0.720000 358.650000 584.600000 358.950000 ;
      RECT 0.000000 353.350000 584.600000 358.650000 ;
      RECT 0.720000 353.050000 584.600000 353.350000 ;
      RECT 0.000000 347.750000 584.600000 353.050000 ;
      RECT 0.720000 347.450000 584.600000 347.750000 ;
      RECT 0.000000 342.150000 584.600000 347.450000 ;
      RECT 0.720000 341.850000 584.600000 342.150000 ;
      RECT 0.000000 336.550000 584.600000 341.850000 ;
      RECT 0.720000 336.250000 584.600000 336.550000 ;
      RECT 0.000000 330.950000 584.600000 336.250000 ;
      RECT 0.720000 330.650000 584.600000 330.950000 ;
      RECT 0.000000 325.350000 584.600000 330.650000 ;
      RECT 0.720000 325.050000 584.600000 325.350000 ;
      RECT 0.000000 319.750000 584.600000 325.050000 ;
      RECT 0.720000 319.450000 584.600000 319.750000 ;
      RECT 0.000000 314.150000 584.600000 319.450000 ;
      RECT 0.720000 313.850000 584.600000 314.150000 ;
      RECT 0.000000 308.550000 584.600000 313.850000 ;
      RECT 0.720000 308.250000 584.600000 308.550000 ;
      RECT 0.000000 302.950000 584.600000 308.250000 ;
      RECT 0.720000 302.650000 584.600000 302.950000 ;
      RECT 0.000000 297.350000 584.600000 302.650000 ;
      RECT 0.720000 297.050000 584.600000 297.350000 ;
      RECT 0.000000 291.750000 584.600000 297.050000 ;
      RECT 0.720000 291.450000 584.600000 291.750000 ;
      RECT 0.000000 286.150000 584.600000 291.450000 ;
      RECT 0.720000 285.850000 584.600000 286.150000 ;
      RECT 0.000000 280.550000 584.600000 285.850000 ;
      RECT 0.720000 280.250000 584.600000 280.550000 ;
      RECT 0.000000 274.950000 584.600000 280.250000 ;
      RECT 0.720000 274.650000 584.600000 274.950000 ;
      RECT 0.000000 269.350000 584.600000 274.650000 ;
      RECT 0.720000 269.050000 584.600000 269.350000 ;
      RECT 0.000000 263.750000 584.600000 269.050000 ;
      RECT 0.720000 263.450000 584.600000 263.750000 ;
      RECT 0.000000 258.150000 584.600000 263.450000 ;
      RECT 0.720000 257.850000 584.600000 258.150000 ;
      RECT 0.000000 252.550000 584.600000 257.850000 ;
      RECT 0.720000 252.250000 584.600000 252.550000 ;
      RECT 0.000000 246.950000 584.600000 252.250000 ;
      RECT 0.720000 246.650000 584.600000 246.950000 ;
      RECT 0.000000 241.350000 584.600000 246.650000 ;
      RECT 0.720000 241.050000 584.600000 241.350000 ;
      RECT 0.000000 235.750000 584.600000 241.050000 ;
      RECT 0.720000 235.450000 584.600000 235.750000 ;
      RECT 0.000000 230.150000 584.600000 235.450000 ;
      RECT 0.720000 229.850000 584.600000 230.150000 ;
      RECT 0.000000 224.550000 584.600000 229.850000 ;
      RECT 0.720000 224.250000 584.600000 224.550000 ;
      RECT 0.000000 218.950000 584.600000 224.250000 ;
      RECT 0.720000 218.650000 584.600000 218.950000 ;
      RECT 0.000000 213.350000 584.600000 218.650000 ;
      RECT 0.720000 213.050000 584.600000 213.350000 ;
      RECT 0.000000 207.750000 584.600000 213.050000 ;
      RECT 0.720000 207.450000 584.600000 207.750000 ;
      RECT 0.000000 202.150000 584.600000 207.450000 ;
      RECT 0.720000 201.850000 584.600000 202.150000 ;
      RECT 0.000000 196.550000 584.600000 201.850000 ;
      RECT 0.720000 196.250000 584.600000 196.550000 ;
      RECT 0.000000 190.750000 584.600000 196.250000 ;
      RECT 0.720000 190.450000 584.600000 190.750000 ;
      RECT 0.000000 185.150000 584.600000 190.450000 ;
      RECT 0.720000 184.850000 584.600000 185.150000 ;
      RECT 0.000000 179.550000 584.600000 184.850000 ;
      RECT 0.720000 179.250000 584.600000 179.550000 ;
      RECT 0.000000 173.950000 584.600000 179.250000 ;
      RECT 0.720000 173.650000 584.600000 173.950000 ;
      RECT 0.000000 168.350000 584.600000 173.650000 ;
      RECT 0.720000 168.050000 584.600000 168.350000 ;
      RECT 0.000000 162.750000 584.600000 168.050000 ;
      RECT 0.720000 162.450000 584.600000 162.750000 ;
      RECT 0.000000 157.150000 584.600000 162.450000 ;
      RECT 0.720000 156.850000 584.600000 157.150000 ;
      RECT 0.000000 151.550000 584.600000 156.850000 ;
      RECT 0.720000 151.250000 584.600000 151.550000 ;
      RECT 0.000000 145.950000 584.600000 151.250000 ;
      RECT 0.720000 145.650000 584.600000 145.950000 ;
      RECT 0.000000 140.350000 584.600000 145.650000 ;
      RECT 0.720000 140.050000 584.600000 140.350000 ;
      RECT 0.000000 134.750000 584.600000 140.050000 ;
      RECT 0.720000 134.450000 584.600000 134.750000 ;
      RECT 0.000000 129.150000 584.600000 134.450000 ;
      RECT 0.720000 128.850000 584.600000 129.150000 ;
      RECT 0.000000 123.550000 584.600000 128.850000 ;
      RECT 0.720000 123.250000 584.600000 123.550000 ;
      RECT 0.000000 117.950000 584.600000 123.250000 ;
      RECT 0.720000 117.650000 584.600000 117.950000 ;
      RECT 0.000000 112.350000 584.600000 117.650000 ;
      RECT 0.720000 112.050000 584.600000 112.350000 ;
      RECT 0.000000 106.750000 584.600000 112.050000 ;
      RECT 0.720000 106.450000 584.600000 106.750000 ;
      RECT 0.000000 101.150000 584.600000 106.450000 ;
      RECT 0.720000 100.850000 584.600000 101.150000 ;
      RECT 0.000000 95.550000 584.600000 100.850000 ;
      RECT 0.720000 95.250000 584.600000 95.550000 ;
      RECT 0.000000 89.950000 584.600000 95.250000 ;
      RECT 0.720000 89.650000 584.600000 89.950000 ;
      RECT 0.000000 84.350000 584.600000 89.650000 ;
      RECT 0.720000 84.050000 584.600000 84.350000 ;
      RECT 0.000000 78.750000 584.600000 84.050000 ;
      RECT 0.720000 78.450000 584.600000 78.750000 ;
      RECT 0.000000 73.150000 584.600000 78.450000 ;
      RECT 0.720000 72.850000 584.600000 73.150000 ;
      RECT 0.000000 67.550000 584.600000 72.850000 ;
      RECT 0.720000 67.250000 584.600000 67.550000 ;
      RECT 0.000000 61.950000 584.600000 67.250000 ;
      RECT 0.720000 61.650000 584.600000 61.950000 ;
      RECT 0.000000 56.350000 584.600000 61.650000 ;
      RECT 0.720000 56.050000 584.600000 56.350000 ;
      RECT 0.000000 50.750000 584.600000 56.050000 ;
      RECT 0.720000 50.450000 584.600000 50.750000 ;
      RECT 0.000000 45.150000 584.600000 50.450000 ;
      RECT 0.720000 44.850000 584.600000 45.150000 ;
      RECT 0.000000 39.550000 584.600000 44.850000 ;
      RECT 0.720000 39.250000 584.600000 39.550000 ;
      RECT 0.000000 33.950000 584.600000 39.250000 ;
      RECT 0.720000 33.650000 584.600000 33.950000 ;
      RECT 0.000000 28.350000 584.600000 33.650000 ;
      RECT 0.720000 28.050000 584.600000 28.350000 ;
      RECT 0.000000 22.750000 584.600000 28.050000 ;
      RECT 0.720000 22.450000 584.600000 22.750000 ;
      RECT 0.000000 17.150000 584.600000 22.450000 ;
      RECT 0.720000 16.850000 584.600000 17.150000 ;
      RECT 0.000000 11.550000 584.600000 16.850000 ;
      RECT 0.720000 11.250000 584.600000 11.550000 ;
      RECT 0.000000 5.950000 584.600000 11.250000 ;
      RECT 0.720000 5.650000 584.600000 5.950000 ;
      RECT 0.000000 0.760000 584.600000 5.650000 ;
      RECT 0.000000 0.350000 0.690000 0.760000 ;
      RECT 581.710000 0.000000 584.290000 0.760000 ;
      RECT 578.710000 0.000000 581.290000 0.760000 ;
      RECT 575.710000 0.000000 578.290000 0.760000 ;
      RECT 572.710000 0.000000 575.290000 0.760000 ;
      RECT 569.910000 0.000000 572.290000 0.760000 ;
      RECT 566.910000 0.000000 569.490000 0.760000 ;
      RECT 563.910000 0.000000 566.490000 0.760000 ;
      RECT 560.910000 0.000000 563.490000 0.760000 ;
      RECT 558.110000 0.000000 560.490000 0.760000 ;
      RECT 555.110000 0.000000 557.690000 0.760000 ;
      RECT 552.110000 0.000000 554.690000 0.760000 ;
      RECT 549.110000 0.000000 551.690000 0.760000 ;
      RECT 546.310000 0.000000 548.690000 0.760000 ;
      RECT 543.310000 0.000000 545.890000 0.760000 ;
      RECT 540.310000 0.000000 542.890000 0.760000 ;
      RECT 537.310000 0.000000 539.890000 0.760000 ;
      RECT 534.510000 0.000000 536.890000 0.760000 ;
      RECT 531.510000 0.000000 534.090000 0.760000 ;
      RECT 528.510000 0.000000 531.090000 0.760000 ;
      RECT 525.510000 0.000000 528.090000 0.760000 ;
      RECT 522.710000 0.000000 525.090000 0.760000 ;
      RECT 519.710000 0.000000 522.290000 0.760000 ;
      RECT 516.710000 0.000000 519.290000 0.760000 ;
      RECT 513.710000 0.000000 516.290000 0.760000 ;
      RECT 510.910000 0.000000 513.290000 0.760000 ;
      RECT 507.910000 0.000000 510.490000 0.760000 ;
      RECT 504.910000 0.000000 507.490000 0.760000 ;
      RECT 501.910000 0.000000 504.490000 0.760000 ;
      RECT 499.110000 0.000000 501.490000 0.760000 ;
      RECT 496.110000 0.000000 498.690000 0.760000 ;
      RECT 493.110000 0.000000 495.690000 0.760000 ;
      RECT 490.110000 0.000000 492.690000 0.760000 ;
      RECT 487.310000 0.000000 489.690000 0.760000 ;
      RECT 484.310000 0.000000 486.890000 0.760000 ;
      RECT 481.310000 0.000000 483.890000 0.760000 ;
      RECT 478.310000 0.000000 480.890000 0.760000 ;
      RECT 475.310000 0.000000 477.890000 0.760000 ;
      RECT 472.510000 0.000000 474.890000 0.760000 ;
      RECT 469.510000 0.000000 472.090000 0.760000 ;
      RECT 466.510000 0.000000 469.090000 0.760000 ;
      RECT 463.510000 0.000000 466.090000 0.760000 ;
      RECT 460.710000 0.000000 463.090000 0.760000 ;
      RECT 457.710000 0.000000 460.290000 0.760000 ;
      RECT 454.710000 0.000000 457.290000 0.760000 ;
      RECT 451.710000 0.000000 454.290000 0.760000 ;
      RECT 448.910000 0.000000 451.290000 0.760000 ;
      RECT 445.910000 0.000000 448.490000 0.760000 ;
      RECT 442.910000 0.000000 445.490000 0.760000 ;
      RECT 439.910000 0.000000 442.490000 0.760000 ;
      RECT 437.110000 0.000000 439.490000 0.760000 ;
      RECT 434.110000 0.000000 436.690000 0.760000 ;
      RECT 431.110000 0.000000 433.690000 0.760000 ;
      RECT 428.110000 0.000000 430.690000 0.760000 ;
      RECT 425.310000 0.000000 427.690000 0.760000 ;
      RECT 422.310000 0.000000 424.890000 0.760000 ;
      RECT 419.310000 0.000000 421.890000 0.760000 ;
      RECT 416.310000 0.000000 418.890000 0.760000 ;
      RECT 413.510000 0.000000 415.890000 0.760000 ;
      RECT 410.510000 0.000000 413.090000 0.760000 ;
      RECT 407.510000 0.000000 410.090000 0.760000 ;
      RECT 404.510000 0.000000 407.090000 0.760000 ;
      RECT 401.710000 0.000000 404.090000 0.760000 ;
      RECT 398.710000 0.000000 401.290000 0.760000 ;
      RECT 395.710000 0.000000 398.290000 0.760000 ;
      RECT 392.710000 0.000000 395.290000 0.760000 ;
      RECT 389.710000 0.000000 392.290000 0.760000 ;
      RECT 386.910000 0.000000 389.290000 0.760000 ;
      RECT 383.910000 0.000000 386.490000 0.760000 ;
      RECT 380.910000 0.000000 383.490000 0.760000 ;
      RECT 377.910000 0.000000 380.490000 0.760000 ;
      RECT 375.110000 0.000000 377.490000 0.760000 ;
      RECT 372.110000 0.000000 374.690000 0.760000 ;
      RECT 369.110000 0.000000 371.690000 0.760000 ;
      RECT 366.110000 0.000000 368.690000 0.760000 ;
      RECT 363.310000 0.000000 365.690000 0.760000 ;
      RECT 360.310000 0.000000 362.890000 0.760000 ;
      RECT 357.310000 0.000000 359.890000 0.760000 ;
      RECT 354.310000 0.000000 356.890000 0.760000 ;
      RECT 351.510000 0.000000 353.890000 0.760000 ;
      RECT 348.510000 0.000000 351.090000 0.760000 ;
      RECT 345.510000 0.000000 348.090000 0.760000 ;
      RECT 342.510000 0.000000 345.090000 0.760000 ;
      RECT 339.710000 0.000000 342.090000 0.760000 ;
      RECT 336.710000 0.000000 339.290000 0.760000 ;
      RECT 333.710000 0.000000 336.290000 0.760000 ;
      RECT 330.710000 0.000000 333.290000 0.760000 ;
      RECT 327.910000 0.000000 330.290000 0.760000 ;
      RECT 324.910000 0.000000 327.490000 0.760000 ;
      RECT 321.910000 0.000000 324.490000 0.760000 ;
      RECT 318.910000 0.000000 321.490000 0.760000 ;
      RECT 316.110000 0.000000 318.490000 0.760000 ;
      RECT 313.110000 0.000000 315.690000 0.760000 ;
      RECT 310.110000 0.000000 312.690000 0.760000 ;
      RECT 307.110000 0.000000 309.690000 0.760000 ;
      RECT 304.310000 0.000000 306.690000 0.760000 ;
      RECT 301.310000 0.000000 303.890000 0.760000 ;
      RECT 298.310000 0.000000 300.890000 0.760000 ;
      RECT 295.310000 0.000000 297.890000 0.760000 ;
      RECT 292.310000 0.000000 294.890000 0.760000 ;
      RECT 289.510000 0.000000 291.890000 0.760000 ;
      RECT 286.510000 0.000000 289.090000 0.760000 ;
      RECT 283.510000 0.000000 286.090000 0.760000 ;
      RECT 280.510000 0.000000 283.090000 0.760000 ;
      RECT 277.710000 0.000000 280.090000 0.760000 ;
      RECT 274.710000 0.000000 277.290000 0.760000 ;
      RECT 271.710000 0.000000 274.290000 0.760000 ;
      RECT 268.710000 0.000000 271.290000 0.760000 ;
      RECT 265.910000 0.000000 268.290000 0.760000 ;
      RECT 262.910000 0.000000 265.490000 0.760000 ;
      RECT 259.910000 0.000000 262.490000 0.760000 ;
      RECT 256.910000 0.000000 259.490000 0.760000 ;
      RECT 254.110000 0.000000 256.490000 0.760000 ;
      RECT 251.110000 0.000000 253.690000 0.760000 ;
      RECT 248.110000 0.000000 250.690000 0.760000 ;
      RECT 245.110000 0.000000 247.690000 0.760000 ;
      RECT 242.310000 0.000000 244.690000 0.760000 ;
      RECT 239.310000 0.000000 241.890000 0.760000 ;
      RECT 236.310000 0.000000 238.890000 0.760000 ;
      RECT 233.310000 0.000000 235.890000 0.760000 ;
      RECT 230.510000 0.000000 232.890000 0.760000 ;
      RECT 227.510000 0.000000 230.090000 0.760000 ;
      RECT 224.510000 0.000000 227.090000 0.760000 ;
      RECT 221.510000 0.000000 224.090000 0.760000 ;
      RECT 218.710000 0.000000 221.090000 0.760000 ;
      RECT 215.710000 0.000000 218.290000 0.760000 ;
      RECT 212.710000 0.000000 215.290000 0.760000 ;
      RECT 209.710000 0.000000 212.290000 0.760000 ;
      RECT 206.910000 0.000000 209.290000 0.760000 ;
      RECT 203.910000 0.000000 206.490000 0.760000 ;
      RECT 200.910000 0.000000 203.490000 0.760000 ;
      RECT 197.910000 0.000000 200.490000 0.760000 ;
      RECT 194.910000 0.000000 197.490000 0.760000 ;
      RECT 192.110000 0.000000 194.490000 0.760000 ;
      RECT 189.110000 0.000000 191.690000 0.760000 ;
      RECT 186.110000 0.000000 188.690000 0.760000 ;
      RECT 183.110000 0.000000 185.690000 0.760000 ;
      RECT 180.310000 0.000000 182.690000 0.760000 ;
      RECT 177.310000 0.000000 179.890000 0.760000 ;
      RECT 174.310000 0.000000 176.890000 0.760000 ;
      RECT 171.310000 0.000000 173.890000 0.760000 ;
      RECT 168.510000 0.000000 170.890000 0.760000 ;
      RECT 165.510000 0.000000 168.090000 0.760000 ;
      RECT 162.510000 0.000000 165.090000 0.760000 ;
      RECT 159.510000 0.000000 162.090000 0.760000 ;
      RECT 156.710000 0.000000 159.090000 0.760000 ;
      RECT 153.710000 0.000000 156.290000 0.760000 ;
      RECT 150.710000 0.000000 153.290000 0.760000 ;
      RECT 147.710000 0.000000 150.290000 0.760000 ;
      RECT 144.910000 0.000000 147.290000 0.760000 ;
      RECT 141.910000 0.000000 144.490000 0.760000 ;
      RECT 138.910000 0.000000 141.490000 0.760000 ;
      RECT 135.910000 0.000000 138.490000 0.760000 ;
      RECT 133.110000 0.000000 135.490000 0.760000 ;
      RECT 130.110000 0.000000 132.690000 0.760000 ;
      RECT 127.110000 0.000000 129.690000 0.760000 ;
      RECT 124.110000 0.000000 126.690000 0.760000 ;
      RECT 121.310000 0.000000 123.690000 0.760000 ;
      RECT 118.310000 0.000000 120.890000 0.760000 ;
      RECT 115.310000 0.000000 117.890000 0.760000 ;
      RECT 112.310000 0.000000 114.890000 0.760000 ;
      RECT 109.510000 0.000000 111.890000 0.760000 ;
      RECT 106.510000 0.000000 109.090000 0.760000 ;
      RECT 103.510000 0.000000 106.090000 0.760000 ;
      RECT 100.510000 0.000000 103.090000 0.760000 ;
      RECT 97.510000 0.000000 100.090000 0.760000 ;
      RECT 94.710000 0.000000 97.090000 0.760000 ;
      RECT 91.710000 0.000000 94.290000 0.760000 ;
      RECT 88.710000 0.000000 91.290000 0.760000 ;
      RECT 85.710000 0.000000 88.290000 0.760000 ;
      RECT 82.910000 0.000000 85.290000 0.760000 ;
      RECT 79.910000 0.000000 82.490000 0.760000 ;
      RECT 76.910000 0.000000 79.490000 0.760000 ;
      RECT 73.910000 0.000000 76.490000 0.760000 ;
      RECT 71.110000 0.000000 73.490000 0.760000 ;
      RECT 68.110000 0.000000 70.690000 0.760000 ;
      RECT 65.110000 0.000000 67.690000 0.760000 ;
      RECT 62.110000 0.000000 64.690000 0.760000 ;
      RECT 59.310000 0.000000 61.690000 0.760000 ;
      RECT 56.310000 0.000000 58.890000 0.760000 ;
      RECT 53.310000 0.000000 55.890000 0.760000 ;
      RECT 50.310000 0.000000 52.890000 0.760000 ;
      RECT 47.510000 0.000000 49.890000 0.760000 ;
      RECT 44.510000 0.000000 47.090000 0.760000 ;
      RECT 41.510000 0.000000 44.090000 0.760000 ;
      RECT 38.510000 0.000000 41.090000 0.760000 ;
      RECT 35.710000 0.000000 38.090000 0.760000 ;
      RECT 32.710000 0.000000 35.290000 0.760000 ;
      RECT 29.710000 0.000000 32.290000 0.760000 ;
      RECT 26.710000 0.000000 29.290000 0.760000 ;
      RECT 23.910000 0.000000 26.290000 0.760000 ;
      RECT 20.910000 0.000000 23.490000 0.760000 ;
      RECT 17.910000 0.000000 20.490000 0.760000 ;
      RECT 14.910000 0.000000 17.490000 0.760000 ;
      RECT 12.110000 0.000000 14.490000 0.760000 ;
      RECT 9.110000 0.000000 11.690000 0.760000 ;
      RECT 6.110000 0.000000 8.690000 0.760000 ;
      RECT 3.110000 0.000000 5.690000 0.760000 ;
      RECT 1.110000 0.000000 2.690000 0.760000 ;
      RECT 0.000000 0.000000 0.690000 0.050000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 584.600000 583.400000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 584.600000 583.400000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 584.600000 583.400000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 584.600000 583.400000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 584.600000 583.400000 ;
  END
END dualcore

END LIBRARY
