##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Thu Mar 23 01:02:28 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO dualcore
  CLASS BLOCK ;
  SIZE 561.600000 BY 558.200000 ;
  FOREIGN dualcore 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 237.700000 0.600000 237.900000 ;
    END
  END clk1
  PIN rst1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 239.300000 0.600000 239.500000 ;
    END
  END rst1
  PIN mem_in_core1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 268.100000 0.600000 268.300000 ;
    END
  END mem_in_core1[31]
  PIN mem_in_core1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 268.900000 0.600000 269.100000 ;
    END
  END mem_in_core1[30]
  PIN mem_in_core1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 269.700000 0.600000 269.900000 ;
    END
  END mem_in_core1[29]
  PIN mem_in_core1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 270.500000 0.600000 270.700000 ;
    END
  END mem_in_core1[28]
  PIN mem_in_core1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 271.300000 0.600000 271.500000 ;
    END
  END mem_in_core1[27]
  PIN mem_in_core1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 272.100000 0.600000 272.300000 ;
    END
  END mem_in_core1[26]
  PIN mem_in_core1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 272.900000 0.600000 273.100000 ;
    END
  END mem_in_core1[25]
  PIN mem_in_core1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 273.700000 0.600000 273.900000 ;
    END
  END mem_in_core1[24]
  PIN mem_in_core1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 274.500000 0.600000 274.700000 ;
    END
  END mem_in_core1[23]
  PIN mem_in_core1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 275.300000 0.600000 275.500000 ;
    END
  END mem_in_core1[22]
  PIN mem_in_core1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 276.100000 0.600000 276.300000 ;
    END
  END mem_in_core1[21]
  PIN mem_in_core1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 276.900000 0.600000 277.100000 ;
    END
  END mem_in_core1[20]
  PIN mem_in_core1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 277.700000 0.600000 277.900000 ;
    END
  END mem_in_core1[19]
  PIN mem_in_core1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 278.500000 0.600000 278.700000 ;
    END
  END mem_in_core1[18]
  PIN mem_in_core1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 279.300000 0.600000 279.500000 ;
    END
  END mem_in_core1[17]
  PIN mem_in_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 280.100000 0.600000 280.300000 ;
    END
  END mem_in_core1[16]
  PIN mem_in_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 280.900000 0.600000 281.100000 ;
    END
  END mem_in_core1[15]
  PIN mem_in_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 281.700000 0.600000 281.900000 ;
    END
  END mem_in_core1[14]
  PIN mem_in_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 282.500000 0.600000 282.700000 ;
    END
  END mem_in_core1[13]
  PIN mem_in_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 283.300000 0.600000 283.500000 ;
    END
  END mem_in_core1[12]
  PIN mem_in_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 284.100000 0.600000 284.300000 ;
    END
  END mem_in_core1[11]
  PIN mem_in_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 284.900000 0.600000 285.100000 ;
    END
  END mem_in_core1[10]
  PIN mem_in_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 285.700000 0.600000 285.900000 ;
    END
  END mem_in_core1[9]
  PIN mem_in_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 286.500000 0.600000 286.700000 ;
    END
  END mem_in_core1[8]
  PIN mem_in_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 287.300000 0.600000 287.500000 ;
    END
  END mem_in_core1[7]
  PIN mem_in_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 288.100000 0.600000 288.300000 ;
    END
  END mem_in_core1[6]
  PIN mem_in_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 288.900000 0.600000 289.100000 ;
    END
  END mem_in_core1[5]
  PIN mem_in_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 289.700000 0.600000 289.900000 ;
    END
  END mem_in_core1[4]
  PIN mem_in_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 290.500000 0.600000 290.700000 ;
    END
  END mem_in_core1[3]
  PIN mem_in_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 291.300000 0.600000 291.500000 ;
    END
  END mem_in_core1[2]
  PIN mem_in_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 292.100000 0.600000 292.300000 ;
    END
  END mem_in_core1[1]
  PIN mem_in_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 292.900000 0.600000 293.100000 ;
    END
  END mem_in_core1[0]
  PIN inst_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 240.900000 0.600000 241.100000 ;
    END
  END inst_core1[16]
  PIN inst_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 241.700000 0.600000 241.900000 ;
    END
  END inst_core1[15]
  PIN inst_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 242.500000 0.600000 242.700000 ;
    END
  END inst_core1[14]
  PIN inst_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 243.300000 0.600000 243.500000 ;
    END
  END inst_core1[13]
  PIN inst_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 244.100000 0.600000 244.300000 ;
    END
  END inst_core1[12]
  PIN inst_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 244.900000 0.600000 245.100000 ;
    END
  END inst_core1[11]
  PIN inst_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 245.700000 0.600000 245.900000 ;
    END
  END inst_core1[10]
  PIN inst_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 246.500000 0.600000 246.700000 ;
    END
  END inst_core1[9]
  PIN inst_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 247.300000 0.600000 247.500000 ;
    END
  END inst_core1[8]
  PIN inst_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 248.100000 0.600000 248.300000 ;
    END
  END inst_core1[7]
  PIN inst_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 248.900000 0.600000 249.100000 ;
    END
  END inst_core1[6]
  PIN inst_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 249.700000 0.600000 249.900000 ;
    END
  END inst_core1[5]
  PIN inst_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 250.500000 0.600000 250.700000 ;
    END
  END inst_core1[4]
  PIN inst_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 251.300000 0.600000 251.500000 ;
    END
  END inst_core1[3]
  PIN inst_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 252.100000 0.600000 252.300000 ;
    END
  END inst_core1[2]
  PIN inst_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 252.900000 0.600000 253.100000 ;
    END
  END inst_core1[1]
  PIN inst_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 253.700000 0.600000 253.900000 ;
    END
  END inst_core1[0]
  PIN out_core1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.800000 0.000000 220.000000 0.600000 ;
    END
  END out_core1[87]
  PIN out_core1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.600000 0.000000 220.800000 0.600000 ;
    END
  END out_core1[86]
  PIN out_core1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 221.400000 0.000000 221.600000 0.600000 ;
    END
  END out_core1[85]
  PIN out_core1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.200000 0.000000 222.400000 0.600000 ;
    END
  END out_core1[84]
  PIN out_core1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.000000 0.000000 223.200000 0.600000 ;
    END
  END out_core1[83]
  PIN out_core1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.800000 0.000000 224.000000 0.600000 ;
    END
  END out_core1[82]
  PIN out_core1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.600000 0.000000 224.800000 0.600000 ;
    END
  END out_core1[81]
  PIN out_core1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 225.400000 0.000000 225.600000 0.600000 ;
    END
  END out_core1[80]
  PIN out_core1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.200000 0.000000 226.400000 0.600000 ;
    END
  END out_core1[79]
  PIN out_core1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.000000 0.000000 227.200000 0.600000 ;
    END
  END out_core1[78]
  PIN out_core1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.800000 0.000000 228.000000 0.600000 ;
    END
  END out_core1[77]
  PIN out_core1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.600000 0.000000 228.800000 0.600000 ;
    END
  END out_core1[76]
  PIN out_core1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.400000 0.000000 229.600000 0.600000 ;
    END
  END out_core1[75]
  PIN out_core1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.200000 0.000000 230.400000 0.600000 ;
    END
  END out_core1[74]
  PIN out_core1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.000000 0.000000 231.200000 0.600000 ;
    END
  END out_core1[73]
  PIN out_core1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.800000 0.000000 232.000000 0.600000 ;
    END
  END out_core1[72]
  PIN out_core1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.600000 0.000000 232.800000 0.600000 ;
    END
  END out_core1[71]
  PIN out_core1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.400000 0.000000 233.600000 0.600000 ;
    END
  END out_core1[70]
  PIN out_core1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.200000 0.000000 234.400000 0.600000 ;
    END
  END out_core1[69]
  PIN out_core1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.000000 0.000000 235.200000 0.600000 ;
    END
  END out_core1[68]
  PIN out_core1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.800000 0.000000 236.000000 0.600000 ;
    END
  END out_core1[67]
  PIN out_core1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 236.600000 0.000000 236.800000 0.600000 ;
    END
  END out_core1[66]
  PIN out_core1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.400000 0.000000 237.600000 0.600000 ;
    END
  END out_core1[65]
  PIN out_core1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.200000 0.000000 238.400000 0.600000 ;
    END
  END out_core1[64]
  PIN out_core1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 239.000000 0.000000 239.200000 0.600000 ;
    END
  END out_core1[63]
  PIN out_core1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 239.800000 0.000000 240.000000 0.600000 ;
    END
  END out_core1[62]
  PIN out_core1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.600000 0.000000 240.800000 0.600000 ;
    END
  END out_core1[61]
  PIN out_core1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.400000 0.000000 241.600000 0.600000 ;
    END
  END out_core1[60]
  PIN out_core1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 242.200000 0.000000 242.400000 0.600000 ;
    END
  END out_core1[59]
  PIN out_core1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.000000 0.000000 243.200000 0.600000 ;
    END
  END out_core1[58]
  PIN out_core1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.800000 0.000000 244.000000 0.600000 ;
    END
  END out_core1[57]
  PIN out_core1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.600000 0.000000 244.800000 0.600000 ;
    END
  END out_core1[56]
  PIN out_core1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.400000 0.000000 245.600000 0.600000 ;
    END
  END out_core1[55]
  PIN out_core1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.200000 0.000000 246.400000 0.600000 ;
    END
  END out_core1[54]
  PIN out_core1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.000000 0.000000 247.200000 0.600000 ;
    END
  END out_core1[53]
  PIN out_core1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.800000 0.000000 248.000000 0.600000 ;
    END
  END out_core1[52]
  PIN out_core1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.600000 0.000000 248.800000 0.600000 ;
    END
  END out_core1[51]
  PIN out_core1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 249.400000 0.000000 249.600000 0.600000 ;
    END
  END out_core1[50]
  PIN out_core1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.200000 0.000000 250.400000 0.600000 ;
    END
  END out_core1[49]
  PIN out_core1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.000000 0.000000 251.200000 0.600000 ;
    END
  END out_core1[48]
  PIN out_core1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.800000 0.000000 252.000000 0.600000 ;
    END
  END out_core1[47]
  PIN out_core1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.600000 0.000000 252.800000 0.600000 ;
    END
  END out_core1[46]
  PIN out_core1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 253.400000 0.000000 253.600000 0.600000 ;
    END
  END out_core1[45]
  PIN out_core1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 254.200000 0.000000 254.400000 0.600000 ;
    END
  END out_core1[44]
  PIN out_core1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.000000 0.000000 255.200000 0.600000 ;
    END
  END out_core1[43]
  PIN out_core1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.800000 0.000000 256.000000 0.600000 ;
    END
  END out_core1[42]
  PIN out_core1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.600000 0.000000 256.800000 0.600000 ;
    END
  END out_core1[41]
  PIN out_core1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 257.400000 0.000000 257.600000 0.600000 ;
    END
  END out_core1[40]
  PIN out_core1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.200000 0.000000 258.400000 0.600000 ;
    END
  END out_core1[39]
  PIN out_core1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.000000 0.000000 259.200000 0.600000 ;
    END
  END out_core1[38]
  PIN out_core1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.800000 0.000000 260.000000 0.600000 ;
    END
  END out_core1[37]
  PIN out_core1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.600000 0.000000 260.800000 0.600000 ;
    END
  END out_core1[36]
  PIN out_core1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.400000 0.000000 261.600000 0.600000 ;
    END
  END out_core1[35]
  PIN out_core1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.200000 0.000000 262.400000 0.600000 ;
    END
  END out_core1[34]
  PIN out_core1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.000000 0.000000 263.200000 0.600000 ;
    END
  END out_core1[33]
  PIN out_core1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.800000 0.000000 264.000000 0.600000 ;
    END
  END out_core1[32]
  PIN out_core1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 264.600000 0.000000 264.800000 0.600000 ;
    END
  END out_core1[31]
  PIN out_core1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.400000 0.000000 265.600000 0.600000 ;
    END
  END out_core1[30]
  PIN out_core1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 266.200000 0.000000 266.400000 0.600000 ;
    END
  END out_core1[29]
  PIN out_core1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.000000 0.000000 267.200000 0.600000 ;
    END
  END out_core1[28]
  PIN out_core1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.800000 0.000000 268.000000 0.600000 ;
    END
  END out_core1[27]
  PIN out_core1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.600000 0.000000 268.800000 0.600000 ;
    END
  END out_core1[26]
  PIN out_core1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 269.400000 0.000000 269.600000 0.600000 ;
    END
  END out_core1[25]
  PIN out_core1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.200000 0.000000 270.400000 0.600000 ;
    END
  END out_core1[24]
  PIN out_core1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.000000 0.000000 271.200000 0.600000 ;
    END
  END out_core1[23]
  PIN out_core1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.800000 0.000000 272.000000 0.600000 ;
    END
  END out_core1[22]
  PIN out_core1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 272.600000 0.000000 272.800000 0.600000 ;
    END
  END out_core1[21]
  PIN out_core1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.400000 0.000000 273.600000 0.600000 ;
    END
  END out_core1[20]
  PIN out_core1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.200000 0.000000 274.400000 0.600000 ;
    END
  END out_core1[19]
  PIN out_core1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.000000 0.000000 275.200000 0.600000 ;
    END
  END out_core1[18]
  PIN out_core1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.800000 0.000000 276.000000 0.600000 ;
    END
  END out_core1[17]
  PIN out_core1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 276.600000 0.000000 276.800000 0.600000 ;
    END
  END out_core1[16]
  PIN out_core1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.400000 0.000000 277.600000 0.600000 ;
    END
  END out_core1[15]
  PIN out_core1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.200000 0.000000 278.400000 0.600000 ;
    END
  END out_core1[14]
  PIN out_core1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.000000 0.000000 279.200000 0.600000 ;
    END
  END out_core1[13]
  PIN out_core1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.800000 0.000000 280.000000 0.600000 ;
    END
  END out_core1[12]
  PIN out_core1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.600000 0.000000 280.800000 0.600000 ;
    END
  END out_core1[11]
  PIN out_core1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.400000 0.000000 281.600000 0.600000 ;
    END
  END out_core1[10]
  PIN out_core1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.200000 0.000000 282.400000 0.600000 ;
    END
  END out_core1[9]
  PIN out_core1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.000000 0.000000 283.200000 0.600000 ;
    END
  END out_core1[8]
  PIN out_core1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.800000 0.000000 284.000000 0.600000 ;
    END
  END out_core1[7]
  PIN out_core1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 284.600000 0.000000 284.800000 0.600000 ;
    END
  END out_core1[6]
  PIN out_core1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.400000 0.000000 285.600000 0.600000 ;
    END
  END out_core1[5]
  PIN out_core1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 286.200000 0.000000 286.400000 0.600000 ;
    END
  END out_core1[4]
  PIN out_core1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.000000 0.000000 287.200000 0.600000 ;
    END
  END out_core1[3]
  PIN out_core1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.800000 0.000000 288.000000 0.600000 ;
    END
  END out_core1[2]
  PIN out_core1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.600000 0.000000 288.800000 0.600000 ;
    END
  END out_core1[1]
  PIN out_core1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.400000 0.000000 289.600000 0.600000 ;
    END
  END out_core1[0]
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 238.500000 0.600000 238.700000 ;
    END
  END clk2
  PIN rst2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 240.100000 0.600000 240.300000 ;
    END
  END rst2
  PIN mem_in_core2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 293.700000 0.600000 293.900000 ;
    END
  END mem_in_core2[31]
  PIN mem_in_core2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 294.500000 0.600000 294.700000 ;
    END
  END mem_in_core2[30]
  PIN mem_in_core2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 295.300000 0.600000 295.500000 ;
    END
  END mem_in_core2[29]
  PIN mem_in_core2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 296.100000 0.600000 296.300000 ;
    END
  END mem_in_core2[28]
  PIN mem_in_core2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 296.900000 0.600000 297.100000 ;
    END
  END mem_in_core2[27]
  PIN mem_in_core2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 297.700000 0.600000 297.900000 ;
    END
  END mem_in_core2[26]
  PIN mem_in_core2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 298.500000 0.600000 298.700000 ;
    END
  END mem_in_core2[25]
  PIN mem_in_core2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 299.300000 0.600000 299.500000 ;
    END
  END mem_in_core2[24]
  PIN mem_in_core2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 300.100000 0.600000 300.300000 ;
    END
  END mem_in_core2[23]
  PIN mem_in_core2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 300.900000 0.600000 301.100000 ;
    END
  END mem_in_core2[22]
  PIN mem_in_core2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 301.700000 0.600000 301.900000 ;
    END
  END mem_in_core2[21]
  PIN mem_in_core2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 302.500000 0.600000 302.700000 ;
    END
  END mem_in_core2[20]
  PIN mem_in_core2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 303.300000 0.600000 303.500000 ;
    END
  END mem_in_core2[19]
  PIN mem_in_core2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.100000 0.600000 304.300000 ;
    END
  END mem_in_core2[18]
  PIN mem_in_core2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.900000 0.600000 305.100000 ;
    END
  END mem_in_core2[17]
  PIN mem_in_core2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 305.700000 0.600000 305.900000 ;
    END
  END mem_in_core2[16]
  PIN mem_in_core2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 306.500000 0.600000 306.700000 ;
    END
  END mem_in_core2[15]
  PIN mem_in_core2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 307.300000 0.600000 307.500000 ;
    END
  END mem_in_core2[14]
  PIN mem_in_core2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 308.100000 0.600000 308.300000 ;
    END
  END mem_in_core2[13]
  PIN mem_in_core2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 308.900000 0.600000 309.100000 ;
    END
  END mem_in_core2[12]
  PIN mem_in_core2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 309.700000 0.600000 309.900000 ;
    END
  END mem_in_core2[11]
  PIN mem_in_core2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 310.500000 0.600000 310.700000 ;
    END
  END mem_in_core2[10]
  PIN mem_in_core2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 311.300000 0.600000 311.500000 ;
    END
  END mem_in_core2[9]
  PIN mem_in_core2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 312.100000 0.600000 312.300000 ;
    END
  END mem_in_core2[8]
  PIN mem_in_core2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 312.900000 0.600000 313.100000 ;
    END
  END mem_in_core2[7]
  PIN mem_in_core2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 313.700000 0.600000 313.900000 ;
    END
  END mem_in_core2[6]
  PIN mem_in_core2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 314.500000 0.600000 314.700000 ;
    END
  END mem_in_core2[5]
  PIN mem_in_core2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 315.300000 0.600000 315.500000 ;
    END
  END mem_in_core2[4]
  PIN mem_in_core2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 316.100000 0.600000 316.300000 ;
    END
  END mem_in_core2[3]
  PIN mem_in_core2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 316.900000 0.600000 317.100000 ;
    END
  END mem_in_core2[2]
  PIN mem_in_core2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 317.700000 0.600000 317.900000 ;
    END
  END mem_in_core2[1]
  PIN mem_in_core2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 318.500000 0.600000 318.700000 ;
    END
  END mem_in_core2[0]
  PIN inst_core2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 254.500000 0.600000 254.700000 ;
    END
  END inst_core2[16]
  PIN inst_core2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 255.300000 0.600000 255.500000 ;
    END
  END inst_core2[15]
  PIN inst_core2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 256.100000 0.600000 256.300000 ;
    END
  END inst_core2[14]
  PIN inst_core2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 256.900000 0.600000 257.100000 ;
    END
  END inst_core2[13]
  PIN inst_core2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 257.700000 0.600000 257.900000 ;
    END
  END inst_core2[12]
  PIN inst_core2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 258.500000 0.600000 258.700000 ;
    END
  END inst_core2[11]
  PIN inst_core2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 259.300000 0.600000 259.500000 ;
    END
  END inst_core2[10]
  PIN inst_core2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 260.100000 0.600000 260.300000 ;
    END
  END inst_core2[9]
  PIN inst_core2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 260.900000 0.600000 261.100000 ;
    END
  END inst_core2[8]
  PIN inst_core2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 261.700000 0.600000 261.900000 ;
    END
  END inst_core2[7]
  PIN inst_core2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 262.500000 0.600000 262.700000 ;
    END
  END inst_core2[6]
  PIN inst_core2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 263.300000 0.600000 263.500000 ;
    END
  END inst_core2[5]
  PIN inst_core2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 264.100000 0.600000 264.300000 ;
    END
  END inst_core2[4]
  PIN inst_core2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 264.900000 0.600000 265.100000 ;
    END
  END inst_core2[3]
  PIN inst_core2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 265.700000 0.600000 265.900000 ;
    END
  END inst_core2[2]
  PIN inst_core2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 266.500000 0.600000 266.700000 ;
    END
  END inst_core2[1]
  PIN inst_core2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 267.300000 0.600000 267.500000 ;
    END
  END inst_core2[0]
  PIN out_core2[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 290.200000 0.000000 290.400000 0.600000 ;
    END
  END out_core2[87]
  PIN out_core2[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.000000 0.000000 291.200000 0.600000 ;
    END
  END out_core2[86]
  PIN out_core2[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.800000 0.000000 292.000000 0.600000 ;
    END
  END out_core2[85]
  PIN out_core2[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 292.600000 0.000000 292.800000 0.600000 ;
    END
  END out_core2[84]
  PIN out_core2[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 293.400000 0.000000 293.600000 0.600000 ;
    END
  END out_core2[83]
  PIN out_core2[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 294.200000 0.000000 294.400000 0.600000 ;
    END
  END out_core2[82]
  PIN out_core2[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.000000 0.000000 295.200000 0.600000 ;
    END
  END out_core2[81]
  PIN out_core2[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.800000 0.000000 296.000000 0.600000 ;
    END
  END out_core2[80]
  PIN out_core2[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 296.600000 0.000000 296.800000 0.600000 ;
    END
  END out_core2[79]
  PIN out_core2[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.400000 0.000000 297.600000 0.600000 ;
    END
  END out_core2[78]
  PIN out_core2[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 298.200000 0.000000 298.400000 0.600000 ;
    END
  END out_core2[77]
  PIN out_core2[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.000000 0.000000 299.200000 0.600000 ;
    END
  END out_core2[76]
  PIN out_core2[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.800000 0.000000 300.000000 0.600000 ;
    END
  END out_core2[75]
  PIN out_core2[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.600000 0.000000 300.800000 0.600000 ;
    END
  END out_core2[74]
  PIN out_core2[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 301.400000 0.000000 301.600000 0.600000 ;
    END
  END out_core2[73]
  PIN out_core2[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.200000 0.000000 302.400000 0.600000 ;
    END
  END out_core2[72]
  PIN out_core2[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.000000 0.000000 303.200000 0.600000 ;
    END
  END out_core2[71]
  PIN out_core2[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.800000 0.000000 304.000000 0.600000 ;
    END
  END out_core2[70]
  PIN out_core2[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 304.600000 0.000000 304.800000 0.600000 ;
    END
  END out_core2[69]
  PIN out_core2[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.400000 0.000000 305.600000 0.600000 ;
    END
  END out_core2[68]
  PIN out_core2[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.200000 0.000000 306.400000 0.600000 ;
    END
  END out_core2[67]
  PIN out_core2[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.000000 0.000000 307.200000 0.600000 ;
    END
  END out_core2[66]
  PIN out_core2[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.800000 0.000000 308.000000 0.600000 ;
    END
  END out_core2[65]
  PIN out_core2[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.600000 0.000000 308.800000 0.600000 ;
    END
  END out_core2[64]
  PIN out_core2[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.400000 0.000000 309.600000 0.600000 ;
    END
  END out_core2[63]
  PIN out_core2[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.200000 0.000000 310.400000 0.600000 ;
    END
  END out_core2[62]
  PIN out_core2[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.000000 0.000000 311.200000 0.600000 ;
    END
  END out_core2[61]
  PIN out_core2[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.800000 0.000000 312.000000 0.600000 ;
    END
  END out_core2[60]
  PIN out_core2[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.600000 0.000000 312.800000 0.600000 ;
    END
  END out_core2[59]
  PIN out_core2[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.400000 0.000000 313.600000 0.600000 ;
    END
  END out_core2[58]
  PIN out_core2[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.200000 0.000000 314.400000 0.600000 ;
    END
  END out_core2[57]
  PIN out_core2[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.000000 0.000000 315.200000 0.600000 ;
    END
  END out_core2[56]
  PIN out_core2[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.800000 0.000000 316.000000 0.600000 ;
    END
  END out_core2[55]
  PIN out_core2[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.600000 0.000000 316.800000 0.600000 ;
    END
  END out_core2[54]
  PIN out_core2[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.400000 0.000000 317.600000 0.600000 ;
    END
  END out_core2[53]
  PIN out_core2[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.200000 0.000000 318.400000 0.600000 ;
    END
  END out_core2[52]
  PIN out_core2[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.000000 0.000000 319.200000 0.600000 ;
    END
  END out_core2[51]
  PIN out_core2[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.800000 0.000000 320.000000 0.600000 ;
    END
  END out_core2[50]
  PIN out_core2[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.600000 0.000000 320.800000 0.600000 ;
    END
  END out_core2[49]
  PIN out_core2[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.400000 0.000000 321.600000 0.600000 ;
    END
  END out_core2[48]
  PIN out_core2[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.200000 0.000000 322.400000 0.600000 ;
    END
  END out_core2[47]
  PIN out_core2[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.000000 0.000000 323.200000 0.600000 ;
    END
  END out_core2[46]
  PIN out_core2[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.800000 0.000000 324.000000 0.600000 ;
    END
  END out_core2[45]
  PIN out_core2[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.600000 0.000000 324.800000 0.600000 ;
    END
  END out_core2[44]
  PIN out_core2[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.400000 0.000000 325.600000 0.600000 ;
    END
  END out_core2[43]
  PIN out_core2[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.200000 0.000000 326.400000 0.600000 ;
    END
  END out_core2[42]
  PIN out_core2[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.000000 0.000000 327.200000 0.600000 ;
    END
  END out_core2[41]
  PIN out_core2[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.800000 0.000000 328.000000 0.600000 ;
    END
  END out_core2[40]
  PIN out_core2[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.600000 0.000000 328.800000 0.600000 ;
    END
  END out_core2[39]
  PIN out_core2[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.400000 0.000000 329.600000 0.600000 ;
    END
  END out_core2[38]
  PIN out_core2[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.200000 0.000000 330.400000 0.600000 ;
    END
  END out_core2[37]
  PIN out_core2[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.000000 0.000000 331.200000 0.600000 ;
    END
  END out_core2[36]
  PIN out_core2[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.800000 0.000000 332.000000 0.600000 ;
    END
  END out_core2[35]
  PIN out_core2[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.600000 0.000000 332.800000 0.600000 ;
    END
  END out_core2[34]
  PIN out_core2[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.400000 0.000000 333.600000 0.600000 ;
    END
  END out_core2[33]
  PIN out_core2[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.200000 0.000000 334.400000 0.600000 ;
    END
  END out_core2[32]
  PIN out_core2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.000000 0.000000 335.200000 0.600000 ;
    END
  END out_core2[31]
  PIN out_core2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.800000 0.000000 336.000000 0.600000 ;
    END
  END out_core2[30]
  PIN out_core2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.600000 0.000000 336.800000 0.600000 ;
    END
  END out_core2[29]
  PIN out_core2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.400000 0.000000 337.600000 0.600000 ;
    END
  END out_core2[28]
  PIN out_core2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.200000 0.000000 338.400000 0.600000 ;
    END
  END out_core2[27]
  PIN out_core2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.000000 0.000000 339.200000 0.600000 ;
    END
  END out_core2[26]
  PIN out_core2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.800000 0.000000 340.000000 0.600000 ;
    END
  END out_core2[25]
  PIN out_core2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.600000 0.000000 340.800000 0.600000 ;
    END
  END out_core2[24]
  PIN out_core2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.400000 0.000000 341.600000 0.600000 ;
    END
  END out_core2[23]
  PIN out_core2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.200000 0.000000 342.400000 0.600000 ;
    END
  END out_core2[22]
  PIN out_core2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.000000 0.000000 343.200000 0.600000 ;
    END
  END out_core2[21]
  PIN out_core2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.800000 0.000000 344.000000 0.600000 ;
    END
  END out_core2[20]
  PIN out_core2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.600000 0.000000 344.800000 0.600000 ;
    END
  END out_core2[19]
  PIN out_core2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.400000 0.000000 345.600000 0.600000 ;
    END
  END out_core2[18]
  PIN out_core2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.200000 0.000000 346.400000 0.600000 ;
    END
  END out_core2[17]
  PIN out_core2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.000000 0.000000 347.200000 0.600000 ;
    END
  END out_core2[16]
  PIN out_core2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.800000 0.000000 348.000000 0.600000 ;
    END
  END out_core2[15]
  PIN out_core2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.600000 0.000000 348.800000 0.600000 ;
    END
  END out_core2[14]
  PIN out_core2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.400000 0.000000 349.600000 0.600000 ;
    END
  END out_core2[13]
  PIN out_core2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.200000 0.000000 350.400000 0.600000 ;
    END
  END out_core2[12]
  PIN out_core2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.000000 0.000000 351.200000 0.600000 ;
    END
  END out_core2[11]
  PIN out_core2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.800000 0.000000 352.000000 0.600000 ;
    END
  END out_core2[10]
  PIN out_core2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.600000 0.000000 352.800000 0.600000 ;
    END
  END out_core2[9]
  PIN out_core2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.400000 0.000000 353.600000 0.600000 ;
    END
  END out_core2[8]
  PIN out_core2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.200000 0.000000 354.400000 0.600000 ;
    END
  END out_core2[7]
  PIN out_core2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.000000 0.000000 355.200000 0.600000 ;
    END
  END out_core2[6]
  PIN out_core2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.800000 0.000000 356.000000 0.600000 ;
    END
  END out_core2[5]
  PIN out_core2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.600000 0.000000 356.800000 0.600000 ;
    END
  END out_core2[4]
  PIN out_core2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.400000 0.000000 357.600000 0.600000 ;
    END
  END out_core2[3]
  PIN out_core2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.200000 0.000000 358.400000 0.600000 ;
    END
  END out_core2[2]
  PIN out_core2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.000000 0.000000 359.200000 0.600000 ;
    END
  END out_core2[1]
  PIN out_core2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.800000 0.000000 360.000000 0.600000 ;
    END
  END out_core2[0]
  PIN s_valid1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 319.300000 0.600000 319.500000 ;
    END
  END s_valid1
  PIN s_valid2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 320.100000 0.600000 320.300000 ;
    END
  END s_valid2
  PIN psum_norm_1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.200000 0.000000 202.400000 0.600000 ;
    END
  END psum_norm_1[10]
  PIN psum_norm_1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.000000 0.000000 203.200000 0.600000 ;
    END
  END psum_norm_1[9]
  PIN psum_norm_1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.800000 0.000000 204.000000 0.600000 ;
    END
  END psum_norm_1[8]
  PIN psum_norm_1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.600000 0.000000 204.800000 0.600000 ;
    END
  END psum_norm_1[7]
  PIN psum_norm_1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.400000 0.000000 205.600000 0.600000 ;
    END
  END psum_norm_1[6]
  PIN psum_norm_1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.200000 0.000000 206.400000 0.600000 ;
    END
  END psum_norm_1[5]
  PIN psum_norm_1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.000000 0.000000 207.200000 0.600000 ;
    END
  END psum_norm_1[4]
  PIN psum_norm_1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.800000 0.000000 208.000000 0.600000 ;
    END
  END psum_norm_1[3]
  PIN psum_norm_1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.600000 0.000000 208.800000 0.600000 ;
    END
  END psum_norm_1[2]
  PIN psum_norm_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.400000 0.000000 209.600000 0.600000 ;
    END
  END psum_norm_1[1]
  PIN psum_norm_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.200000 0.000000 210.400000 0.600000 ;
    END
  END psum_norm_1[0]
  PIN psum_norm_2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.000000 0.000000 211.200000 0.600000 ;
    END
  END psum_norm_2[10]
  PIN psum_norm_2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.800000 0.000000 212.000000 0.600000 ;
    END
  END psum_norm_2[9]
  PIN psum_norm_2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.600000 0.000000 212.800000 0.600000 ;
    END
  END psum_norm_2[8]
  PIN psum_norm_2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.400000 0.000000 213.600000 0.600000 ;
    END
  END psum_norm_2[7]
  PIN psum_norm_2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.200000 0.000000 214.400000 0.600000 ;
    END
  END psum_norm_2[6]
  PIN psum_norm_2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.000000 0.000000 215.200000 0.600000 ;
    END
  END psum_norm_2[5]
  PIN psum_norm_2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.800000 0.000000 216.000000 0.600000 ;
    END
  END psum_norm_2[4]
  PIN psum_norm_2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.600000 0.000000 216.800000 0.600000 ;
    END
  END psum_norm_2[3]
  PIN psum_norm_2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.400000 0.000000 217.600000 0.600000 ;
    END
  END psum_norm_2[2]
  PIN psum_norm_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.200000 0.000000 218.400000 0.600000 ;
    END
  END psum_norm_2[1]
  PIN psum_norm_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.000000 0.000000 219.200000 0.600000 ;
    END
  END psum_norm_2[0]
  PIN norm_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.400000 0.000000 201.600000 0.600000 ;
    END
  END norm_valid
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 561.600000 558.200000 ;
    LAYER M2 ;
      RECT 0.000000 0.700000 561.600000 558.200000 ;
      RECT 360.100000 0.000000 561.600000 0.700000 ;
      RECT 359.300000 0.000000 359.700000 0.700000 ;
      RECT 358.500000 0.000000 358.900000 0.700000 ;
      RECT 357.700000 0.000000 358.100000 0.700000 ;
      RECT 356.900000 0.000000 357.300000 0.700000 ;
      RECT 356.100000 0.000000 356.500000 0.700000 ;
      RECT 355.300000 0.000000 355.700000 0.700000 ;
      RECT 354.500000 0.000000 354.900000 0.700000 ;
      RECT 353.700000 0.000000 354.100000 0.700000 ;
      RECT 352.900000 0.000000 353.300000 0.700000 ;
      RECT 352.100000 0.000000 352.500000 0.700000 ;
      RECT 351.300000 0.000000 351.700000 0.700000 ;
      RECT 350.500000 0.000000 350.900000 0.700000 ;
      RECT 349.700000 0.000000 350.100000 0.700000 ;
      RECT 348.900000 0.000000 349.300000 0.700000 ;
      RECT 348.100000 0.000000 348.500000 0.700000 ;
      RECT 347.300000 0.000000 347.700000 0.700000 ;
      RECT 346.500000 0.000000 346.900000 0.700000 ;
      RECT 345.700000 0.000000 346.100000 0.700000 ;
      RECT 344.900000 0.000000 345.300000 0.700000 ;
      RECT 344.100000 0.000000 344.500000 0.700000 ;
      RECT 343.300000 0.000000 343.700000 0.700000 ;
      RECT 342.500000 0.000000 342.900000 0.700000 ;
      RECT 341.700000 0.000000 342.100000 0.700000 ;
      RECT 340.900000 0.000000 341.300000 0.700000 ;
      RECT 340.100000 0.000000 340.500000 0.700000 ;
      RECT 339.300000 0.000000 339.700000 0.700000 ;
      RECT 338.500000 0.000000 338.900000 0.700000 ;
      RECT 337.700000 0.000000 338.100000 0.700000 ;
      RECT 336.900000 0.000000 337.300000 0.700000 ;
      RECT 336.100000 0.000000 336.500000 0.700000 ;
      RECT 335.300000 0.000000 335.700000 0.700000 ;
      RECT 334.500000 0.000000 334.900000 0.700000 ;
      RECT 333.700000 0.000000 334.100000 0.700000 ;
      RECT 332.900000 0.000000 333.300000 0.700000 ;
      RECT 332.100000 0.000000 332.500000 0.700000 ;
      RECT 331.300000 0.000000 331.700000 0.700000 ;
      RECT 330.500000 0.000000 330.900000 0.700000 ;
      RECT 329.700000 0.000000 330.100000 0.700000 ;
      RECT 328.900000 0.000000 329.300000 0.700000 ;
      RECT 328.100000 0.000000 328.500000 0.700000 ;
      RECT 327.300000 0.000000 327.700000 0.700000 ;
      RECT 326.500000 0.000000 326.900000 0.700000 ;
      RECT 325.700000 0.000000 326.100000 0.700000 ;
      RECT 324.900000 0.000000 325.300000 0.700000 ;
      RECT 324.100000 0.000000 324.500000 0.700000 ;
      RECT 323.300000 0.000000 323.700000 0.700000 ;
      RECT 322.500000 0.000000 322.900000 0.700000 ;
      RECT 321.700000 0.000000 322.100000 0.700000 ;
      RECT 320.900000 0.000000 321.300000 0.700000 ;
      RECT 320.100000 0.000000 320.500000 0.700000 ;
      RECT 319.300000 0.000000 319.700000 0.700000 ;
      RECT 318.500000 0.000000 318.900000 0.700000 ;
      RECT 317.700000 0.000000 318.100000 0.700000 ;
      RECT 316.900000 0.000000 317.300000 0.700000 ;
      RECT 316.100000 0.000000 316.500000 0.700000 ;
      RECT 315.300000 0.000000 315.700000 0.700000 ;
      RECT 314.500000 0.000000 314.900000 0.700000 ;
      RECT 313.700000 0.000000 314.100000 0.700000 ;
      RECT 312.900000 0.000000 313.300000 0.700000 ;
      RECT 312.100000 0.000000 312.500000 0.700000 ;
      RECT 311.300000 0.000000 311.700000 0.700000 ;
      RECT 310.500000 0.000000 310.900000 0.700000 ;
      RECT 309.700000 0.000000 310.100000 0.700000 ;
      RECT 308.900000 0.000000 309.300000 0.700000 ;
      RECT 308.100000 0.000000 308.500000 0.700000 ;
      RECT 307.300000 0.000000 307.700000 0.700000 ;
      RECT 306.500000 0.000000 306.900000 0.700000 ;
      RECT 305.700000 0.000000 306.100000 0.700000 ;
      RECT 304.900000 0.000000 305.300000 0.700000 ;
      RECT 304.100000 0.000000 304.500000 0.700000 ;
      RECT 303.300000 0.000000 303.700000 0.700000 ;
      RECT 302.500000 0.000000 302.900000 0.700000 ;
      RECT 301.700000 0.000000 302.100000 0.700000 ;
      RECT 300.900000 0.000000 301.300000 0.700000 ;
      RECT 300.100000 0.000000 300.500000 0.700000 ;
      RECT 299.300000 0.000000 299.700000 0.700000 ;
      RECT 298.500000 0.000000 298.900000 0.700000 ;
      RECT 297.700000 0.000000 298.100000 0.700000 ;
      RECT 296.900000 0.000000 297.300000 0.700000 ;
      RECT 296.100000 0.000000 296.500000 0.700000 ;
      RECT 295.300000 0.000000 295.700000 0.700000 ;
      RECT 294.500000 0.000000 294.900000 0.700000 ;
      RECT 293.700000 0.000000 294.100000 0.700000 ;
      RECT 292.900000 0.000000 293.300000 0.700000 ;
      RECT 292.100000 0.000000 292.500000 0.700000 ;
      RECT 291.300000 0.000000 291.700000 0.700000 ;
      RECT 290.500000 0.000000 290.900000 0.700000 ;
      RECT 289.700000 0.000000 290.100000 0.700000 ;
      RECT 288.900000 0.000000 289.300000 0.700000 ;
      RECT 288.100000 0.000000 288.500000 0.700000 ;
      RECT 287.300000 0.000000 287.700000 0.700000 ;
      RECT 286.500000 0.000000 286.900000 0.700000 ;
      RECT 285.700000 0.000000 286.100000 0.700000 ;
      RECT 284.900000 0.000000 285.300000 0.700000 ;
      RECT 284.100000 0.000000 284.500000 0.700000 ;
      RECT 283.300000 0.000000 283.700000 0.700000 ;
      RECT 282.500000 0.000000 282.900000 0.700000 ;
      RECT 281.700000 0.000000 282.100000 0.700000 ;
      RECT 280.900000 0.000000 281.300000 0.700000 ;
      RECT 280.100000 0.000000 280.500000 0.700000 ;
      RECT 279.300000 0.000000 279.700000 0.700000 ;
      RECT 278.500000 0.000000 278.900000 0.700000 ;
      RECT 277.700000 0.000000 278.100000 0.700000 ;
      RECT 276.900000 0.000000 277.300000 0.700000 ;
      RECT 276.100000 0.000000 276.500000 0.700000 ;
      RECT 275.300000 0.000000 275.700000 0.700000 ;
      RECT 274.500000 0.000000 274.900000 0.700000 ;
      RECT 273.700000 0.000000 274.100000 0.700000 ;
      RECT 272.900000 0.000000 273.300000 0.700000 ;
      RECT 272.100000 0.000000 272.500000 0.700000 ;
      RECT 271.300000 0.000000 271.700000 0.700000 ;
      RECT 270.500000 0.000000 270.900000 0.700000 ;
      RECT 269.700000 0.000000 270.100000 0.700000 ;
      RECT 268.900000 0.000000 269.300000 0.700000 ;
      RECT 268.100000 0.000000 268.500000 0.700000 ;
      RECT 267.300000 0.000000 267.700000 0.700000 ;
      RECT 266.500000 0.000000 266.900000 0.700000 ;
      RECT 265.700000 0.000000 266.100000 0.700000 ;
      RECT 264.900000 0.000000 265.300000 0.700000 ;
      RECT 264.100000 0.000000 264.500000 0.700000 ;
      RECT 263.300000 0.000000 263.700000 0.700000 ;
      RECT 262.500000 0.000000 262.900000 0.700000 ;
      RECT 261.700000 0.000000 262.100000 0.700000 ;
      RECT 260.900000 0.000000 261.300000 0.700000 ;
      RECT 260.100000 0.000000 260.500000 0.700000 ;
      RECT 259.300000 0.000000 259.700000 0.700000 ;
      RECT 258.500000 0.000000 258.900000 0.700000 ;
      RECT 257.700000 0.000000 258.100000 0.700000 ;
      RECT 256.900000 0.000000 257.300000 0.700000 ;
      RECT 256.100000 0.000000 256.500000 0.700000 ;
      RECT 255.300000 0.000000 255.700000 0.700000 ;
      RECT 254.500000 0.000000 254.900000 0.700000 ;
      RECT 253.700000 0.000000 254.100000 0.700000 ;
      RECT 252.900000 0.000000 253.300000 0.700000 ;
      RECT 252.100000 0.000000 252.500000 0.700000 ;
      RECT 251.300000 0.000000 251.700000 0.700000 ;
      RECT 250.500000 0.000000 250.900000 0.700000 ;
      RECT 249.700000 0.000000 250.100000 0.700000 ;
      RECT 248.900000 0.000000 249.300000 0.700000 ;
      RECT 248.100000 0.000000 248.500000 0.700000 ;
      RECT 247.300000 0.000000 247.700000 0.700000 ;
      RECT 246.500000 0.000000 246.900000 0.700000 ;
      RECT 245.700000 0.000000 246.100000 0.700000 ;
      RECT 244.900000 0.000000 245.300000 0.700000 ;
      RECT 244.100000 0.000000 244.500000 0.700000 ;
      RECT 243.300000 0.000000 243.700000 0.700000 ;
      RECT 242.500000 0.000000 242.900000 0.700000 ;
      RECT 241.700000 0.000000 242.100000 0.700000 ;
      RECT 240.900000 0.000000 241.300000 0.700000 ;
      RECT 240.100000 0.000000 240.500000 0.700000 ;
      RECT 239.300000 0.000000 239.700000 0.700000 ;
      RECT 238.500000 0.000000 238.900000 0.700000 ;
      RECT 237.700000 0.000000 238.100000 0.700000 ;
      RECT 236.900000 0.000000 237.300000 0.700000 ;
      RECT 236.100000 0.000000 236.500000 0.700000 ;
      RECT 235.300000 0.000000 235.700000 0.700000 ;
      RECT 234.500000 0.000000 234.900000 0.700000 ;
      RECT 233.700000 0.000000 234.100000 0.700000 ;
      RECT 232.900000 0.000000 233.300000 0.700000 ;
      RECT 232.100000 0.000000 232.500000 0.700000 ;
      RECT 231.300000 0.000000 231.700000 0.700000 ;
      RECT 230.500000 0.000000 230.900000 0.700000 ;
      RECT 229.700000 0.000000 230.100000 0.700000 ;
      RECT 228.900000 0.000000 229.300000 0.700000 ;
      RECT 228.100000 0.000000 228.500000 0.700000 ;
      RECT 227.300000 0.000000 227.700000 0.700000 ;
      RECT 226.500000 0.000000 226.900000 0.700000 ;
      RECT 225.700000 0.000000 226.100000 0.700000 ;
      RECT 224.900000 0.000000 225.300000 0.700000 ;
      RECT 224.100000 0.000000 224.500000 0.700000 ;
      RECT 223.300000 0.000000 223.700000 0.700000 ;
      RECT 222.500000 0.000000 222.900000 0.700000 ;
      RECT 221.700000 0.000000 222.100000 0.700000 ;
      RECT 220.900000 0.000000 221.300000 0.700000 ;
      RECT 220.100000 0.000000 220.500000 0.700000 ;
      RECT 219.300000 0.000000 219.700000 0.700000 ;
      RECT 218.500000 0.000000 218.900000 0.700000 ;
      RECT 217.700000 0.000000 218.100000 0.700000 ;
      RECT 216.900000 0.000000 217.300000 0.700000 ;
      RECT 216.100000 0.000000 216.500000 0.700000 ;
      RECT 215.300000 0.000000 215.700000 0.700000 ;
      RECT 214.500000 0.000000 214.900000 0.700000 ;
      RECT 213.700000 0.000000 214.100000 0.700000 ;
      RECT 212.900000 0.000000 213.300000 0.700000 ;
      RECT 212.100000 0.000000 212.500000 0.700000 ;
      RECT 211.300000 0.000000 211.700000 0.700000 ;
      RECT 210.500000 0.000000 210.900000 0.700000 ;
      RECT 209.700000 0.000000 210.100000 0.700000 ;
      RECT 208.900000 0.000000 209.300000 0.700000 ;
      RECT 208.100000 0.000000 208.500000 0.700000 ;
      RECT 207.300000 0.000000 207.700000 0.700000 ;
      RECT 206.500000 0.000000 206.900000 0.700000 ;
      RECT 205.700000 0.000000 206.100000 0.700000 ;
      RECT 204.900000 0.000000 205.300000 0.700000 ;
      RECT 204.100000 0.000000 204.500000 0.700000 ;
      RECT 203.300000 0.000000 203.700000 0.700000 ;
      RECT 202.500000 0.000000 202.900000 0.700000 ;
      RECT 201.700000 0.000000 202.100000 0.700000 ;
      RECT 0.000000 0.000000 201.300000 0.700000 ;
    LAYER M3 ;
      RECT 0.000000 320.400000 561.600000 558.200000 ;
      RECT 0.700000 320.000000 561.600000 320.400000 ;
      RECT 0.000000 319.600000 561.600000 320.000000 ;
      RECT 0.700000 319.200000 561.600000 319.600000 ;
      RECT 0.000000 318.800000 561.600000 319.200000 ;
      RECT 0.700000 318.400000 561.600000 318.800000 ;
      RECT 0.000000 318.000000 561.600000 318.400000 ;
      RECT 0.700000 317.600000 561.600000 318.000000 ;
      RECT 0.000000 317.200000 561.600000 317.600000 ;
      RECT 0.700000 316.800000 561.600000 317.200000 ;
      RECT 0.000000 316.400000 561.600000 316.800000 ;
      RECT 0.700000 316.000000 561.600000 316.400000 ;
      RECT 0.000000 315.600000 561.600000 316.000000 ;
      RECT 0.700000 315.200000 561.600000 315.600000 ;
      RECT 0.000000 314.800000 561.600000 315.200000 ;
      RECT 0.700000 314.400000 561.600000 314.800000 ;
      RECT 0.000000 314.000000 561.600000 314.400000 ;
      RECT 0.700000 313.600000 561.600000 314.000000 ;
      RECT 0.000000 313.200000 561.600000 313.600000 ;
      RECT 0.700000 312.800000 561.600000 313.200000 ;
      RECT 0.000000 312.400000 561.600000 312.800000 ;
      RECT 0.700000 312.000000 561.600000 312.400000 ;
      RECT 0.000000 311.600000 561.600000 312.000000 ;
      RECT 0.700000 311.200000 561.600000 311.600000 ;
      RECT 0.000000 310.800000 561.600000 311.200000 ;
      RECT 0.700000 310.400000 561.600000 310.800000 ;
      RECT 0.000000 310.000000 561.600000 310.400000 ;
      RECT 0.700000 309.600000 561.600000 310.000000 ;
      RECT 0.000000 309.200000 561.600000 309.600000 ;
      RECT 0.700000 308.800000 561.600000 309.200000 ;
      RECT 0.000000 308.400000 561.600000 308.800000 ;
      RECT 0.700000 308.000000 561.600000 308.400000 ;
      RECT 0.000000 307.600000 561.600000 308.000000 ;
      RECT 0.700000 307.200000 561.600000 307.600000 ;
      RECT 0.000000 306.800000 561.600000 307.200000 ;
      RECT 0.700000 306.400000 561.600000 306.800000 ;
      RECT 0.000000 306.000000 561.600000 306.400000 ;
      RECT 0.700000 305.600000 561.600000 306.000000 ;
      RECT 0.000000 305.200000 561.600000 305.600000 ;
      RECT 0.700000 304.800000 561.600000 305.200000 ;
      RECT 0.000000 304.400000 561.600000 304.800000 ;
      RECT 0.700000 304.000000 561.600000 304.400000 ;
      RECT 0.000000 303.600000 561.600000 304.000000 ;
      RECT 0.700000 303.200000 561.600000 303.600000 ;
      RECT 0.000000 302.800000 561.600000 303.200000 ;
      RECT 0.700000 302.400000 561.600000 302.800000 ;
      RECT 0.000000 302.000000 561.600000 302.400000 ;
      RECT 0.700000 301.600000 561.600000 302.000000 ;
      RECT 0.000000 301.200000 561.600000 301.600000 ;
      RECT 0.700000 300.800000 561.600000 301.200000 ;
      RECT 0.000000 300.400000 561.600000 300.800000 ;
      RECT 0.700000 300.000000 561.600000 300.400000 ;
      RECT 0.000000 299.600000 561.600000 300.000000 ;
      RECT 0.700000 299.200000 561.600000 299.600000 ;
      RECT 0.000000 298.800000 561.600000 299.200000 ;
      RECT 0.700000 298.400000 561.600000 298.800000 ;
      RECT 0.000000 298.000000 561.600000 298.400000 ;
      RECT 0.700000 297.600000 561.600000 298.000000 ;
      RECT 0.000000 297.200000 561.600000 297.600000 ;
      RECT 0.700000 296.800000 561.600000 297.200000 ;
      RECT 0.000000 296.400000 561.600000 296.800000 ;
      RECT 0.700000 296.000000 561.600000 296.400000 ;
      RECT 0.000000 295.600000 561.600000 296.000000 ;
      RECT 0.700000 295.200000 561.600000 295.600000 ;
      RECT 0.000000 294.800000 561.600000 295.200000 ;
      RECT 0.700000 294.400000 561.600000 294.800000 ;
      RECT 0.000000 294.000000 561.600000 294.400000 ;
      RECT 0.700000 293.600000 561.600000 294.000000 ;
      RECT 0.000000 293.200000 561.600000 293.600000 ;
      RECT 0.700000 292.800000 561.600000 293.200000 ;
      RECT 0.000000 292.400000 561.600000 292.800000 ;
      RECT 0.700000 292.000000 561.600000 292.400000 ;
      RECT 0.000000 291.600000 561.600000 292.000000 ;
      RECT 0.700000 291.200000 561.600000 291.600000 ;
      RECT 0.000000 290.800000 561.600000 291.200000 ;
      RECT 0.700000 290.400000 561.600000 290.800000 ;
      RECT 0.000000 290.000000 561.600000 290.400000 ;
      RECT 0.700000 289.600000 561.600000 290.000000 ;
      RECT 0.000000 289.200000 561.600000 289.600000 ;
      RECT 0.700000 288.800000 561.600000 289.200000 ;
      RECT 0.000000 288.400000 561.600000 288.800000 ;
      RECT 0.700000 288.000000 561.600000 288.400000 ;
      RECT 0.000000 287.600000 561.600000 288.000000 ;
      RECT 0.700000 287.200000 561.600000 287.600000 ;
      RECT 0.000000 286.800000 561.600000 287.200000 ;
      RECT 0.700000 286.400000 561.600000 286.800000 ;
      RECT 0.000000 286.000000 561.600000 286.400000 ;
      RECT 0.700000 285.600000 561.600000 286.000000 ;
      RECT 0.000000 285.200000 561.600000 285.600000 ;
      RECT 0.700000 284.800000 561.600000 285.200000 ;
      RECT 0.000000 284.400000 561.600000 284.800000 ;
      RECT 0.700000 284.000000 561.600000 284.400000 ;
      RECT 0.000000 283.600000 561.600000 284.000000 ;
      RECT 0.700000 283.200000 561.600000 283.600000 ;
      RECT 0.000000 282.800000 561.600000 283.200000 ;
      RECT 0.700000 282.400000 561.600000 282.800000 ;
      RECT 0.000000 282.000000 561.600000 282.400000 ;
      RECT 0.700000 281.600000 561.600000 282.000000 ;
      RECT 0.000000 281.200000 561.600000 281.600000 ;
      RECT 0.700000 280.800000 561.600000 281.200000 ;
      RECT 0.000000 280.400000 561.600000 280.800000 ;
      RECT 0.700000 280.000000 561.600000 280.400000 ;
      RECT 0.000000 279.600000 561.600000 280.000000 ;
      RECT 0.700000 279.200000 561.600000 279.600000 ;
      RECT 0.000000 278.800000 561.600000 279.200000 ;
      RECT 0.700000 278.400000 561.600000 278.800000 ;
      RECT 0.000000 278.000000 561.600000 278.400000 ;
      RECT 0.700000 277.600000 561.600000 278.000000 ;
      RECT 0.000000 277.200000 561.600000 277.600000 ;
      RECT 0.700000 276.800000 561.600000 277.200000 ;
      RECT 0.000000 276.400000 561.600000 276.800000 ;
      RECT 0.700000 276.000000 561.600000 276.400000 ;
      RECT 0.000000 275.600000 561.600000 276.000000 ;
      RECT 0.700000 275.200000 561.600000 275.600000 ;
      RECT 0.000000 274.800000 561.600000 275.200000 ;
      RECT 0.700000 274.400000 561.600000 274.800000 ;
      RECT 0.000000 274.000000 561.600000 274.400000 ;
      RECT 0.700000 273.600000 561.600000 274.000000 ;
      RECT 0.000000 273.200000 561.600000 273.600000 ;
      RECT 0.700000 272.800000 561.600000 273.200000 ;
      RECT 0.000000 272.400000 561.600000 272.800000 ;
      RECT 0.700000 272.000000 561.600000 272.400000 ;
      RECT 0.000000 271.600000 561.600000 272.000000 ;
      RECT 0.700000 271.200000 561.600000 271.600000 ;
      RECT 0.000000 270.800000 561.600000 271.200000 ;
      RECT 0.700000 270.400000 561.600000 270.800000 ;
      RECT 0.000000 270.000000 561.600000 270.400000 ;
      RECT 0.700000 269.600000 561.600000 270.000000 ;
      RECT 0.000000 269.200000 561.600000 269.600000 ;
      RECT 0.700000 268.800000 561.600000 269.200000 ;
      RECT 0.000000 268.400000 561.600000 268.800000 ;
      RECT 0.700000 268.000000 561.600000 268.400000 ;
      RECT 0.000000 267.600000 561.600000 268.000000 ;
      RECT 0.700000 267.200000 561.600000 267.600000 ;
      RECT 0.000000 266.800000 561.600000 267.200000 ;
      RECT 0.700000 266.400000 561.600000 266.800000 ;
      RECT 0.000000 266.000000 561.600000 266.400000 ;
      RECT 0.700000 265.600000 561.600000 266.000000 ;
      RECT 0.000000 265.200000 561.600000 265.600000 ;
      RECT 0.700000 264.800000 561.600000 265.200000 ;
      RECT 0.000000 264.400000 561.600000 264.800000 ;
      RECT 0.700000 264.000000 561.600000 264.400000 ;
      RECT 0.000000 263.600000 561.600000 264.000000 ;
      RECT 0.700000 263.200000 561.600000 263.600000 ;
      RECT 0.000000 262.800000 561.600000 263.200000 ;
      RECT 0.700000 262.400000 561.600000 262.800000 ;
      RECT 0.000000 262.000000 561.600000 262.400000 ;
      RECT 0.700000 261.600000 561.600000 262.000000 ;
      RECT 0.000000 261.200000 561.600000 261.600000 ;
      RECT 0.700000 260.800000 561.600000 261.200000 ;
      RECT 0.000000 260.400000 561.600000 260.800000 ;
      RECT 0.700000 260.000000 561.600000 260.400000 ;
      RECT 0.000000 259.600000 561.600000 260.000000 ;
      RECT 0.700000 259.200000 561.600000 259.600000 ;
      RECT 0.000000 258.800000 561.600000 259.200000 ;
      RECT 0.700000 258.400000 561.600000 258.800000 ;
      RECT 0.000000 258.000000 561.600000 258.400000 ;
      RECT 0.700000 257.600000 561.600000 258.000000 ;
      RECT 0.000000 257.200000 561.600000 257.600000 ;
      RECT 0.700000 256.800000 561.600000 257.200000 ;
      RECT 0.000000 256.400000 561.600000 256.800000 ;
      RECT 0.700000 256.000000 561.600000 256.400000 ;
      RECT 0.000000 255.600000 561.600000 256.000000 ;
      RECT 0.700000 255.200000 561.600000 255.600000 ;
      RECT 0.000000 254.800000 561.600000 255.200000 ;
      RECT 0.700000 254.400000 561.600000 254.800000 ;
      RECT 0.000000 254.000000 561.600000 254.400000 ;
      RECT 0.700000 253.600000 561.600000 254.000000 ;
      RECT 0.000000 253.200000 561.600000 253.600000 ;
      RECT 0.700000 252.800000 561.600000 253.200000 ;
      RECT 0.000000 252.400000 561.600000 252.800000 ;
      RECT 0.700000 252.000000 561.600000 252.400000 ;
      RECT 0.000000 251.600000 561.600000 252.000000 ;
      RECT 0.700000 251.200000 561.600000 251.600000 ;
      RECT 0.000000 250.800000 561.600000 251.200000 ;
      RECT 0.700000 250.400000 561.600000 250.800000 ;
      RECT 0.000000 250.000000 561.600000 250.400000 ;
      RECT 0.700000 249.600000 561.600000 250.000000 ;
      RECT 0.000000 249.200000 561.600000 249.600000 ;
      RECT 0.700000 248.800000 561.600000 249.200000 ;
      RECT 0.000000 248.400000 561.600000 248.800000 ;
      RECT 0.700000 248.000000 561.600000 248.400000 ;
      RECT 0.000000 247.600000 561.600000 248.000000 ;
      RECT 0.700000 247.200000 561.600000 247.600000 ;
      RECT 0.000000 246.800000 561.600000 247.200000 ;
      RECT 0.700000 246.400000 561.600000 246.800000 ;
      RECT 0.000000 246.000000 561.600000 246.400000 ;
      RECT 0.700000 245.600000 561.600000 246.000000 ;
      RECT 0.000000 245.200000 561.600000 245.600000 ;
      RECT 0.700000 244.800000 561.600000 245.200000 ;
      RECT 0.000000 244.400000 561.600000 244.800000 ;
      RECT 0.700000 244.000000 561.600000 244.400000 ;
      RECT 0.000000 243.600000 561.600000 244.000000 ;
      RECT 0.700000 243.200000 561.600000 243.600000 ;
      RECT 0.000000 242.800000 561.600000 243.200000 ;
      RECT 0.700000 242.400000 561.600000 242.800000 ;
      RECT 0.000000 242.000000 561.600000 242.400000 ;
      RECT 0.700000 241.600000 561.600000 242.000000 ;
      RECT 0.000000 241.200000 561.600000 241.600000 ;
      RECT 0.700000 240.800000 561.600000 241.200000 ;
      RECT 0.000000 240.400000 561.600000 240.800000 ;
      RECT 0.700000 240.000000 561.600000 240.400000 ;
      RECT 0.000000 239.600000 561.600000 240.000000 ;
      RECT 0.700000 239.200000 561.600000 239.600000 ;
      RECT 0.000000 238.800000 561.600000 239.200000 ;
      RECT 0.700000 238.400000 561.600000 238.800000 ;
      RECT 0.000000 238.000000 561.600000 238.400000 ;
      RECT 0.700000 237.600000 561.600000 238.000000 ;
      RECT 0.000000 0.000000 561.600000 237.600000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 561.600000 558.200000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 561.600000 558.200000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 561.600000 558.200000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 561.600000 558.200000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 561.600000 558.200000 ;
  END
END dualcore

END LIBRARY
