##
## LEF for PtnCells ;
<<<<<<< HEAD
## created by Innovus v19.17-s077_1 on Thu Mar 23 08:44:44 2023
=======
## created by Innovus v19.17-s077_1 on Thu Mar 23 12:36:34 2023
>>>>>>> aed9910e876bdd4365d7eb9a7bdff198e5814b9b
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO dualcore
  CLASS BLOCK ;
  SIZE 568.000000 BY 565.400000 ;
  FOREIGN dualcore 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 460.500000 0.600000 460.700000 ;
    END
  END clk1
  PIN rst1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 457.300000 0.600000 457.500000 ;
    END
  END rst1
  PIN mem_in_core1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 428.500000 0.600000 428.700000 ;
    END
  END mem_in_core1[31]
  PIN mem_in_core1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 427.700000 0.600000 427.900000 ;
    END
  END mem_in_core1[30]
  PIN mem_in_core1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 426.900000 0.600000 427.100000 ;
    END
  END mem_in_core1[29]
  PIN mem_in_core1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 426.100000 0.600000 426.300000 ;
    END
  END mem_in_core1[28]
  PIN mem_in_core1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 425.300000 0.600000 425.500000 ;
    END
  END mem_in_core1[27]
  PIN mem_in_core1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 424.500000 0.600000 424.700000 ;
    END
  END mem_in_core1[26]
  PIN mem_in_core1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 423.700000 0.600000 423.900000 ;
    END
  END mem_in_core1[25]
  PIN mem_in_core1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 422.900000 0.600000 423.100000 ;
    END
  END mem_in_core1[24]
  PIN mem_in_core1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 422.100000 0.600000 422.300000 ;
    END
  END mem_in_core1[23]
  PIN mem_in_core1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 421.300000 0.600000 421.500000 ;
    END
  END mem_in_core1[22]
  PIN mem_in_core1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 420.500000 0.600000 420.700000 ;
    END
  END mem_in_core1[21]
  PIN mem_in_core1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 419.700000 0.600000 419.900000 ;
    END
  END mem_in_core1[20]
  PIN mem_in_core1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 418.900000 0.600000 419.100000 ;
    END
  END mem_in_core1[19]
  PIN mem_in_core1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 418.100000 0.600000 418.300000 ;
    END
  END mem_in_core1[18]
  PIN mem_in_core1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 417.300000 0.600000 417.500000 ;
    END
  END mem_in_core1[17]
  PIN mem_in_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 416.500000 0.600000 416.700000 ;
    END
  END mem_in_core1[16]
  PIN mem_in_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 415.700000 0.600000 415.900000 ;
    END
  END mem_in_core1[15]
  PIN mem_in_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 414.900000 0.600000 415.100000 ;
    END
  END mem_in_core1[14]
  PIN mem_in_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 414.100000 0.600000 414.300000 ;
    END
  END mem_in_core1[13]
  PIN mem_in_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 413.300000 0.600000 413.500000 ;
    END
  END mem_in_core1[12]
  PIN mem_in_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 412.500000 0.600000 412.700000 ;
    END
  END mem_in_core1[11]
  PIN mem_in_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 411.700000 0.600000 411.900000 ;
    END
  END mem_in_core1[10]
  PIN mem_in_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 410.900000 0.600000 411.100000 ;
    END
  END mem_in_core1[9]
  PIN mem_in_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 410.100000 0.600000 410.300000 ;
    END
  END mem_in_core1[8]
  PIN mem_in_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 409.300000 0.600000 409.500000 ;
    END
  END mem_in_core1[7]
  PIN mem_in_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 408.500000 0.600000 408.700000 ;
    END
  END mem_in_core1[6]
  PIN mem_in_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 407.700000 0.600000 407.900000 ;
    END
  END mem_in_core1[5]
  PIN mem_in_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 406.900000 0.600000 407.100000 ;
    END
  END mem_in_core1[4]
  PIN mem_in_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 406.100000 0.600000 406.300000 ;
    END
  END mem_in_core1[3]
  PIN mem_in_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 405.300000 0.600000 405.500000 ;
    END
  END mem_in_core1[2]
  PIN mem_in_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 404.500000 0.600000 404.700000 ;
    END
  END mem_in_core1[1]
  PIN mem_in_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 403.700000 0.600000 403.900000 ;
    END
  END mem_in_core1[0]
  PIN inst_core1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 455.700000 0.600000 455.900000 ;
    END
  END inst_core1[16]
  PIN inst_core1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 454.900000 0.600000 455.100000 ;
    END
  END inst_core1[15]
  PIN inst_core1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 454.100000 0.600000 454.300000 ;
    END
  END inst_core1[14]
  PIN inst_core1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 453.300000 0.600000 453.500000 ;
    END
  END inst_core1[13]
  PIN inst_core1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 452.500000 0.600000 452.700000 ;
    END
  END inst_core1[12]
  PIN inst_core1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 451.700000 0.600000 451.900000 ;
    END
  END inst_core1[11]
  PIN inst_core1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 450.900000 0.600000 451.100000 ;
    END
  END inst_core1[10]
  PIN inst_core1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 450.100000 0.600000 450.300000 ;
    END
  END inst_core1[9]
  PIN inst_core1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 449.300000 0.600000 449.500000 ;
    END
  END inst_core1[8]
  PIN inst_core1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 448.500000 0.600000 448.700000 ;
    END
  END inst_core1[7]
  PIN inst_core1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 447.700000 0.600000 447.900000 ;
    END
  END inst_core1[6]
  PIN inst_core1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 446.900000 0.600000 447.100000 ;
    END
  END inst_core1[5]
  PIN inst_core1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 446.100000 0.600000 446.300000 ;
    END
  END inst_core1[4]
  PIN inst_core1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 445.300000 0.600000 445.500000 ;
    END
  END inst_core1[3]
  PIN inst_core1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 444.500000 0.600000 444.700000 ;
    END
  END inst_core1[2]
  PIN inst_core1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 443.700000 0.600000 443.900000 ;
    END
  END inst_core1[1]
  PIN inst_core1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 442.900000 0.600000 443.100000 ;
    END
  END inst_core1[0]
  PIN out_core1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.400000 0.000000 440.600000 0.600000 ;
    END
  END out_core1[87]
  PIN out_core1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.600000 0.000000 439.800000 0.600000 ;
    END
  END out_core1[86]
  PIN out_core1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.800000 0.000000 439.000000 0.600000 ;
    END
  END out_core1[85]
  PIN out_core1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.000000 0.000000 438.200000 0.600000 ;
    END
  END out_core1[84]
  PIN out_core1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 437.200000 0.000000 437.400000 0.600000 ;
    END
  END out_core1[83]
  PIN out_core1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.400000 0.000000 436.600000 0.600000 ;
    END
  END out_core1[82]
  PIN out_core1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.600000 0.000000 435.800000 0.600000 ;
    END
  END out_core1[81]
  PIN out_core1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.800000 0.000000 435.000000 0.600000 ;
    END
  END out_core1[80]
  PIN out_core1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.000000 0.000000 434.200000 0.600000 ;
    END
  END out_core1[79]
  PIN out_core1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.200000 0.000000 433.400000 0.600000 ;
    END
  END out_core1[78]
  PIN out_core1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.400000 0.000000 432.600000 0.600000 ;
    END
  END out_core1[77]
  PIN out_core1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.600000 0.000000 431.800000 0.600000 ;
    END
  END out_core1[76]
  PIN out_core1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.800000 0.000000 431.000000 0.600000 ;
    END
  END out_core1[75]
  PIN out_core1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.000000 0.000000 430.200000 0.600000 ;
    END
  END out_core1[74]
  PIN out_core1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 429.200000 0.000000 429.400000 0.600000 ;
    END
  END out_core1[73]
  PIN out_core1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.400000 0.000000 428.600000 0.600000 ;
    END
  END out_core1[72]
  PIN out_core1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.600000 0.000000 427.800000 0.600000 ;
    END
  END out_core1[71]
  PIN out_core1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.800000 0.000000 427.000000 0.600000 ;
    END
  END out_core1[70]
  PIN out_core1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.000000 0.000000 426.200000 0.600000 ;
    END
  END out_core1[69]
  PIN out_core1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.200000 0.000000 425.400000 0.600000 ;
    END
  END out_core1[68]
  PIN out_core1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.400000 0.000000 424.600000 0.600000 ;
    END
  END out_core1[67]
  PIN out_core1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.600000 0.000000 423.800000 0.600000 ;
    END
  END out_core1[66]
  PIN out_core1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.800000 0.000000 423.000000 0.600000 ;
    END
  END out_core1[65]
  PIN out_core1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.000000 0.000000 422.200000 0.600000 ;
    END
  END out_core1[64]
  PIN out_core1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 421.200000 0.000000 421.400000 0.600000 ;
    END
  END out_core1[63]
  PIN out_core1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.400000 0.000000 420.600000 0.600000 ;
    END
  END out_core1[62]
  PIN out_core1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.600000 0.000000 419.800000 0.600000 ;
    END
  END out_core1[61]
  PIN out_core1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.800000 0.000000 419.000000 0.600000 ;
    END
  END out_core1[60]
  PIN out_core1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.000000 0.000000 418.200000 0.600000 ;
    END
  END out_core1[59]
  PIN out_core1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.200000 0.000000 417.400000 0.600000 ;
    END
  END out_core1[58]
  PIN out_core1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 416.400000 0.000000 416.600000 0.600000 ;
    END
  END out_core1[57]
  PIN out_core1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.600000 0.000000 415.800000 0.600000 ;
    END
  END out_core1[56]
  PIN out_core1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.800000 0.000000 415.000000 0.600000 ;
    END
  END out_core1[55]
  PIN out_core1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.000000 0.000000 414.200000 0.600000 ;
    END
  END out_core1[54]
  PIN out_core1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 413.200000 0.000000 413.400000 0.600000 ;
    END
  END out_core1[53]
  PIN out_core1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.400000 0.000000 412.600000 0.600000 ;
    END
  END out_core1[52]
  PIN out_core1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.600000 0.000000 411.800000 0.600000 ;
    END
  END out_core1[51]
  PIN out_core1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.800000 0.000000 411.000000 0.600000 ;
    END
  END out_core1[50]
  PIN out_core1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.000000 0.000000 410.200000 0.600000 ;
    END
  END out_core1[49]
  PIN out_core1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 409.200000 0.000000 409.400000 0.600000 ;
    END
  END out_core1[48]
  PIN out_core1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.400000 0.000000 408.600000 0.600000 ;
    END
  END out_core1[47]
  PIN out_core1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.600000 0.000000 407.800000 0.600000 ;
    END
  END out_core1[46]
  PIN out_core1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.800000 0.000000 407.000000 0.600000 ;
    END
  END out_core1[45]
  PIN out_core1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.000000 0.000000 406.200000 0.600000 ;
    END
  END out_core1[44]
  PIN out_core1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.200000 0.000000 405.400000 0.600000 ;
    END
  END out_core1[43]
  PIN out_core1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.400000 0.000000 404.600000 0.600000 ;
    END
  END out_core1[42]
  PIN out_core1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.600000 0.000000 403.800000 0.600000 ;
    END
  END out_core1[41]
  PIN out_core1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.800000 0.000000 403.000000 0.600000 ;
    END
  END out_core1[40]
  PIN out_core1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.000000 0.000000 402.200000 0.600000 ;
    END
  END out_core1[39]
  PIN out_core1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 401.200000 0.000000 401.400000 0.600000 ;
    END
  END out_core1[38]
  PIN out_core1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.400000 0.000000 400.600000 0.600000 ;
    END
  END out_core1[37]
  PIN out_core1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.600000 0.000000 399.800000 0.600000 ;
    END
  END out_core1[36]
  PIN out_core1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.800000 0.000000 399.000000 0.600000 ;
    END
  END out_core1[35]
  PIN out_core1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.000000 0.000000 398.200000 0.600000 ;
    END
  END out_core1[34]
  PIN out_core1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.200000 0.000000 397.400000 0.600000 ;
    END
  END out_core1[33]
  PIN out_core1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.400000 0.000000 396.600000 0.600000 ;
    END
  END out_core1[32]
  PIN out_core1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.600000 0.000000 395.800000 0.600000 ;
    END
  END out_core1[31]
  PIN out_core1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.800000 0.000000 395.000000 0.600000 ;
    END
  END out_core1[30]
  PIN out_core1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.000000 0.000000 394.200000 0.600000 ;
    END
  END out_core1[29]
  PIN out_core1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 393.200000 0.000000 393.400000 0.600000 ;
    END
  END out_core1[28]
  PIN out_core1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.400000 0.000000 392.600000 0.600000 ;
    END
  END out_core1[27]
  PIN out_core1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.600000 0.000000 391.800000 0.600000 ;
    END
  END out_core1[26]
  PIN out_core1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.800000 0.000000 391.000000 0.600000 ;
    END
  END out_core1[25]
  PIN out_core1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.000000 0.000000 390.200000 0.600000 ;
    END
  END out_core1[24]
  PIN out_core1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.200000 0.000000 389.400000 0.600000 ;
    END
  END out_core1[23]
  PIN out_core1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.400000 0.000000 388.600000 0.600000 ;
    END
  END out_core1[22]
  PIN out_core1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.600000 0.000000 387.800000 0.600000 ;
    END
  END out_core1[21]
  PIN out_core1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.800000 0.000000 387.000000 0.600000 ;
    END
  END out_core1[20]
  PIN out_core1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.000000 0.000000 386.200000 0.600000 ;
    END
  END out_core1[19]
  PIN out_core1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.200000 0.000000 385.400000 0.600000 ;
    END
  END out_core1[18]
  PIN out_core1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.400000 0.000000 384.600000 0.600000 ;
    END
  END out_core1[17]
  PIN out_core1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.600000 0.000000 383.800000 0.600000 ;
    END
  END out_core1[16]
  PIN out_core1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.800000 0.000000 383.000000 0.600000 ;
    END
  END out_core1[15]
  PIN out_core1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.000000 0.000000 382.200000 0.600000 ;
    END
  END out_core1[14]
  PIN out_core1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.200000 0.000000 381.400000 0.600000 ;
    END
  END out_core1[13]
  PIN out_core1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.400000 0.000000 380.600000 0.600000 ;
    END
  END out_core1[12]
  PIN out_core1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.600000 0.000000 379.800000 0.600000 ;
    END
  END out_core1[11]
  PIN out_core1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.800000 0.000000 379.000000 0.600000 ;
    END
  END out_core1[10]
  PIN out_core1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.000000 0.000000 378.200000 0.600000 ;
    END
  END out_core1[9]
  PIN out_core1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 377.200000 0.000000 377.400000 0.600000 ;
    END
  END out_core1[8]
  PIN out_core1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.400000 0.000000 376.600000 0.600000 ;
    END
  END out_core1[7]
  PIN out_core1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.600000 0.000000 375.800000 0.600000 ;
    END
  END out_core1[6]
  PIN out_core1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.800000 0.000000 375.000000 0.600000 ;
    END
  END out_core1[5]
  PIN out_core1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.000000 0.000000 374.200000 0.600000 ;
    END
  END out_core1[4]
  PIN out_core1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.200000 0.000000 373.400000 0.600000 ;
    END
  END out_core1[3]
  PIN out_core1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.400000 0.000000 372.600000 0.600000 ;
    END
  END out_core1[2]
  PIN out_core1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.600000 0.000000 371.800000 0.600000 ;
    END
  END out_core1[1]
  PIN out_core1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.800000 0.000000 371.000000 0.600000 ;
    END
  END out_core1[0]
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 459.700000 0.600000 459.900000 ;
    END
  END clk2
  PIN rst2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 456.500000 0.600000 456.700000 ;
    END
  END rst2
  PIN mem_in_core2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 402.900000 0.600000 403.100000 ;
    END
  END mem_in_core2[31]
  PIN mem_in_core2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 402.100000 0.600000 402.300000 ;
    END
  END mem_in_core2[30]
  PIN mem_in_core2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 401.300000 0.600000 401.500000 ;
    END
  END mem_in_core2[29]
  PIN mem_in_core2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 400.500000 0.600000 400.700000 ;
    END
  END mem_in_core2[28]
  PIN mem_in_core2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 399.700000 0.600000 399.900000 ;
    END
  END mem_in_core2[27]
  PIN mem_in_core2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 398.900000 0.600000 399.100000 ;
    END
  END mem_in_core2[26]
  PIN mem_in_core2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 398.100000 0.600000 398.300000 ;
    END
  END mem_in_core2[25]
  PIN mem_in_core2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 397.300000 0.600000 397.500000 ;
    END
  END mem_in_core2[24]
  PIN mem_in_core2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 396.500000 0.600000 396.700000 ;
    END
  END mem_in_core2[23]
  PIN mem_in_core2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 395.700000 0.600000 395.900000 ;
    END
  END mem_in_core2[22]
  PIN mem_in_core2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 394.900000 0.600000 395.100000 ;
    END
  END mem_in_core2[21]
  PIN mem_in_core2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 394.100000 0.600000 394.300000 ;
    END
  END mem_in_core2[20]
  PIN mem_in_core2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 393.300000 0.600000 393.500000 ;
    END
  END mem_in_core2[19]
  PIN mem_in_core2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 392.500000 0.600000 392.700000 ;
    END
  END mem_in_core2[18]
  PIN mem_in_core2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 391.700000 0.600000 391.900000 ;
    END
  END mem_in_core2[17]
  PIN mem_in_core2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 390.900000 0.600000 391.100000 ;
    END
  END mem_in_core2[16]
  PIN mem_in_core2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 390.100000 0.600000 390.300000 ;
    END
  END mem_in_core2[15]
  PIN mem_in_core2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 389.300000 0.600000 389.500000 ;
    END
  END mem_in_core2[14]
  PIN mem_in_core2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 388.500000 0.600000 388.700000 ;
    END
  END mem_in_core2[13]
  PIN mem_in_core2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 387.700000 0.600000 387.900000 ;
    END
  END mem_in_core2[12]
  PIN mem_in_core2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 386.900000 0.600000 387.100000 ;
    END
  END mem_in_core2[11]
  PIN mem_in_core2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 386.100000 0.600000 386.300000 ;
    END
  END mem_in_core2[10]
  PIN mem_in_core2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 385.300000 0.600000 385.500000 ;
    END
  END mem_in_core2[9]
  PIN mem_in_core2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 384.500000 0.600000 384.700000 ;
    END
  END mem_in_core2[8]
  PIN mem_in_core2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 383.700000 0.600000 383.900000 ;
    END
  END mem_in_core2[7]
  PIN mem_in_core2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 382.900000 0.600000 383.100000 ;
    END
  END mem_in_core2[6]
  PIN mem_in_core2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 382.100000 0.600000 382.300000 ;
    END
  END mem_in_core2[5]
  PIN mem_in_core2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 381.300000 0.600000 381.500000 ;
    END
  END mem_in_core2[4]
  PIN mem_in_core2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 380.500000 0.600000 380.700000 ;
    END
  END mem_in_core2[3]
  PIN mem_in_core2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 379.700000 0.600000 379.900000 ;
    END
  END mem_in_core2[2]
  PIN mem_in_core2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 378.900000 0.600000 379.100000 ;
    END
  END mem_in_core2[1]
  PIN mem_in_core2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 378.100000 0.600000 378.300000 ;
    END
  END mem_in_core2[0]
  PIN inst_core2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 442.100000 0.600000 442.300000 ;
    END
  END inst_core2[16]
  PIN inst_core2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 441.300000 0.600000 441.500000 ;
    END
  END inst_core2[15]
  PIN inst_core2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 440.500000 0.600000 440.700000 ;
    END
  END inst_core2[14]
  PIN inst_core2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 439.700000 0.600000 439.900000 ;
    END
  END inst_core2[13]
  PIN inst_core2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 438.900000 0.600000 439.100000 ;
    END
  END inst_core2[12]
  PIN inst_core2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 438.100000 0.600000 438.300000 ;
    END
  END inst_core2[11]
  PIN inst_core2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 437.300000 0.600000 437.500000 ;
    END
  END inst_core2[10]
  PIN inst_core2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 436.500000 0.600000 436.700000 ;
    END
  END inst_core2[9]
  PIN inst_core2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 435.700000 0.600000 435.900000 ;
    END
  END inst_core2[8]
  PIN inst_core2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 434.900000 0.600000 435.100000 ;
    END
  END inst_core2[7]
  PIN inst_core2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 434.100000 0.600000 434.300000 ;
    END
  END inst_core2[6]
  PIN inst_core2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 433.300000 0.600000 433.500000 ;
    END
  END inst_core2[5]
  PIN inst_core2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 432.500000 0.600000 432.700000 ;
    END
  END inst_core2[4]
  PIN inst_core2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 431.700000 0.600000 431.900000 ;
    END
  END inst_core2[3]
  PIN inst_core2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 430.900000 0.600000 431.100000 ;
    END
  END inst_core2[2]
  PIN inst_core2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 430.100000 0.600000 430.300000 ;
    END
  END inst_core2[1]
  PIN inst_core2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 429.300000 0.600000 429.500000 ;
    END
  END inst_core2[0]
  PIN out_core2[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.000000 0.000000 370.200000 0.600000 ;
    END
  END out_core2[87]
  PIN out_core2[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.200000 0.000000 369.400000 0.600000 ;
    END
  END out_core2[86]
  PIN out_core2[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.400000 0.000000 368.600000 0.600000 ;
    END
  END out_core2[85]
  PIN out_core2[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.600000 0.000000 367.800000 0.600000 ;
    END
  END out_core2[84]
  PIN out_core2[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.800000 0.000000 367.000000 0.600000 ;
    END
  END out_core2[83]
  PIN out_core2[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.000000 0.000000 366.200000 0.600000 ;
    END
  END out_core2[82]
  PIN out_core2[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.200000 0.000000 365.400000 0.600000 ;
    END
  END out_core2[81]
  PIN out_core2[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.400000 0.000000 364.600000 0.600000 ;
    END
  END out_core2[80]
  PIN out_core2[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.600000 0.000000 363.800000 0.600000 ;
    END
  END out_core2[79]
  PIN out_core2[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.800000 0.000000 363.000000 0.600000 ;
    END
  END out_core2[78]
  PIN out_core2[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.000000 0.000000 362.200000 0.600000 ;
    END
  END out_core2[77]
  PIN out_core2[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.200000 0.000000 361.400000 0.600000 ;
    END
  END out_core2[76]
  PIN out_core2[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.400000 0.000000 360.600000 0.600000 ;
    END
  END out_core2[75]
  PIN out_core2[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.600000 0.000000 359.800000 0.600000 ;
    END
  END out_core2[74]
  PIN out_core2[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.800000 0.000000 359.000000 0.600000 ;
    END
  END out_core2[73]
  PIN out_core2[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.000000 0.000000 358.200000 0.600000 ;
    END
  END out_core2[72]
  PIN out_core2[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.200000 0.000000 357.400000 0.600000 ;
    END
  END out_core2[71]
  PIN out_core2[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.400000 0.000000 356.600000 0.600000 ;
    END
  END out_core2[70]
  PIN out_core2[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.600000 0.000000 355.800000 0.600000 ;
    END
  END out_core2[69]
  PIN out_core2[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.800000 0.000000 355.000000 0.600000 ;
    END
  END out_core2[68]
  PIN out_core2[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.000000 0.000000 354.200000 0.600000 ;
    END
  END out_core2[67]
  PIN out_core2[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.200000 0.000000 353.400000 0.600000 ;
    END
  END out_core2[66]
  PIN out_core2[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.400000 0.000000 352.600000 0.600000 ;
    END
  END out_core2[65]
  PIN out_core2[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.600000 0.000000 351.800000 0.600000 ;
    END
  END out_core2[64]
  PIN out_core2[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.800000 0.000000 351.000000 0.600000 ;
    END
  END out_core2[63]
  PIN out_core2[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.000000 0.000000 350.200000 0.600000 ;
    END
  END out_core2[62]
  PIN out_core2[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.200000 0.000000 349.400000 0.600000 ;
    END
  END out_core2[61]
  PIN out_core2[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.400000 0.000000 348.600000 0.600000 ;
    END
  END out_core2[60]
  PIN out_core2[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.600000 0.000000 347.800000 0.600000 ;
    END
  END out_core2[59]
  PIN out_core2[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.800000 0.000000 347.000000 0.600000 ;
    END
  END out_core2[58]
  PIN out_core2[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.000000 0.000000 346.200000 0.600000 ;
    END
  END out_core2[57]
  PIN out_core2[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.200000 0.000000 345.400000 0.600000 ;
    END
  END out_core2[56]
  PIN out_core2[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.400000 0.000000 344.600000 0.600000 ;
    END
  END out_core2[55]
  PIN out_core2[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.600000 0.000000 343.800000 0.600000 ;
    END
  END out_core2[54]
  PIN out_core2[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.800000 0.000000 343.000000 0.600000 ;
    END
  END out_core2[53]
  PIN out_core2[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.000000 0.000000 342.200000 0.600000 ;
    END
  END out_core2[52]
  PIN out_core2[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.200000 0.000000 341.400000 0.600000 ;
    END
  END out_core2[51]
  PIN out_core2[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.400000 0.000000 340.600000 0.600000 ;
    END
  END out_core2[50]
  PIN out_core2[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.600000 0.000000 339.800000 0.600000 ;
    END
  END out_core2[49]
  PIN out_core2[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.800000 0.000000 339.000000 0.600000 ;
    END
  END out_core2[48]
  PIN out_core2[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.000000 0.000000 338.200000 0.600000 ;
    END
  END out_core2[47]
  PIN out_core2[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.200000 0.000000 337.400000 0.600000 ;
    END
  END out_core2[46]
  PIN out_core2[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.400000 0.000000 336.600000 0.600000 ;
    END
  END out_core2[45]
  PIN out_core2[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.600000 0.000000 335.800000 0.600000 ;
    END
  END out_core2[44]
  PIN out_core2[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.800000 0.000000 335.000000 0.600000 ;
    END
  END out_core2[43]
  PIN out_core2[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.000000 0.000000 334.200000 0.600000 ;
    END
  END out_core2[42]
  PIN out_core2[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.200000 0.000000 333.400000 0.600000 ;
    END
  END out_core2[41]
  PIN out_core2[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.400000 0.000000 332.600000 0.600000 ;
    END
  END out_core2[40]
  PIN out_core2[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.600000 0.000000 331.800000 0.600000 ;
    END
  END out_core2[39]
  PIN out_core2[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.800000 0.000000 331.000000 0.600000 ;
    END
  END out_core2[38]
  PIN out_core2[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.000000 0.000000 330.200000 0.600000 ;
    END
  END out_core2[37]
  PIN out_core2[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.200000 0.000000 329.400000 0.600000 ;
    END
  END out_core2[36]
  PIN out_core2[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.400000 0.000000 328.600000 0.600000 ;
    END
  END out_core2[35]
  PIN out_core2[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.600000 0.000000 327.800000 0.600000 ;
    END
  END out_core2[34]
  PIN out_core2[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.800000 0.000000 327.000000 0.600000 ;
    END
  END out_core2[33]
  PIN out_core2[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.000000 0.000000 326.200000 0.600000 ;
    END
  END out_core2[32]
  PIN out_core2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.200000 0.000000 325.400000 0.600000 ;
    END
  END out_core2[31]
  PIN out_core2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.400000 0.000000 324.600000 0.600000 ;
    END
  END out_core2[30]
  PIN out_core2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.600000 0.000000 323.800000 0.600000 ;
    END
  END out_core2[29]
  PIN out_core2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.800000 0.000000 323.000000 0.600000 ;
    END
  END out_core2[28]
  PIN out_core2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.000000 0.000000 322.200000 0.600000 ;
    END
  END out_core2[27]
  PIN out_core2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.200000 0.000000 321.400000 0.600000 ;
    END
  END out_core2[26]
  PIN out_core2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.400000 0.000000 320.600000 0.600000 ;
    END
  END out_core2[25]
  PIN out_core2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.600000 0.000000 319.800000 0.600000 ;
    END
  END out_core2[24]
  PIN out_core2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.800000 0.000000 319.000000 0.600000 ;
    END
  END out_core2[23]
  PIN out_core2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.000000 0.000000 318.200000 0.600000 ;
    END
  END out_core2[22]
  PIN out_core2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.200000 0.000000 317.400000 0.600000 ;
    END
  END out_core2[21]
  PIN out_core2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.400000 0.000000 316.600000 0.600000 ;
    END
  END out_core2[20]
  PIN out_core2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.600000 0.000000 315.800000 0.600000 ;
    END
  END out_core2[19]
  PIN out_core2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.800000 0.000000 315.000000 0.600000 ;
    END
  END out_core2[18]
  PIN out_core2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.000000 0.000000 314.200000 0.600000 ;
    END
  END out_core2[17]
  PIN out_core2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.200000 0.000000 313.400000 0.600000 ;
    END
  END out_core2[16]
  PIN out_core2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.400000 0.000000 312.600000 0.600000 ;
    END
  END out_core2[15]
  PIN out_core2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.600000 0.000000 311.800000 0.600000 ;
    END
  END out_core2[14]
  PIN out_core2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.800000 0.000000 311.000000 0.600000 ;
    END
  END out_core2[13]
  PIN out_core2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.000000 0.000000 310.200000 0.600000 ;
    END
  END out_core2[12]
  PIN out_core2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.200000 0.000000 309.400000 0.600000 ;
    END
  END out_core2[11]
  PIN out_core2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.400000 0.000000 308.600000 0.600000 ;
    END
  END out_core2[10]
  PIN out_core2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.600000 0.000000 307.800000 0.600000 ;
    END
  END out_core2[9]
  PIN out_core2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.800000 0.000000 307.000000 0.600000 ;
    END
  END out_core2[8]
  PIN out_core2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.000000 0.000000 306.200000 0.600000 ;
    END
  END out_core2[7]
  PIN out_core2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.200000 0.000000 305.400000 0.600000 ;
    END
  END out_core2[6]
  PIN out_core2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 304.400000 0.000000 304.600000 0.600000 ;
    END
  END out_core2[5]
  PIN out_core2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.600000 0.000000 303.800000 0.600000 ;
    END
  END out_core2[4]
  PIN out_core2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.800000 0.000000 303.000000 0.600000 ;
    END
  END out_core2[3]
  PIN out_core2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.000000 0.000000 302.200000 0.600000 ;
    END
  END out_core2[2]
  PIN out_core2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 301.200000 0.000000 301.400000 0.600000 ;
    END
  END out_core2[1]
  PIN out_core2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.400000 0.000000 300.600000 0.600000 ;
    END
  END out_core2[0]
  PIN core_gate1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 458.900000 0.600000 459.100000 ;
    END
  END core_gate1
  PIN core_gate2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 458.100000 0.600000 458.300000 ;
    END
  END core_gate2
  PIN s_valid1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 460.400000 0.000000 460.600000 0.600000 ;
    END
  END s_valid1
  PIN s_valid2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 459.600000 0.000000 459.800000 0.600000 ;
    END
  END s_valid2
  PIN psum_norm_1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 458.000000 0.000000 458.200000 0.600000 ;
    END
  END psum_norm_1[10]
  PIN psum_norm_1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.200000 0.000000 457.400000 0.600000 ;
    END
  END psum_norm_1[9]
  PIN psum_norm_1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.400000 0.000000 456.600000 0.600000 ;
    END
  END psum_norm_1[8]
  PIN psum_norm_1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.600000 0.000000 455.800000 0.600000 ;
    END
  END psum_norm_1[7]
  PIN psum_norm_1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.800000 0.000000 455.000000 0.600000 ;
    END
  END psum_norm_1[6]
  PIN psum_norm_1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.000000 0.000000 454.200000 0.600000 ;
    END
  END psum_norm_1[5]
  PIN psum_norm_1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 453.200000 0.000000 453.400000 0.600000 ;
    END
  END psum_norm_1[4]
  PIN psum_norm_1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.400000 0.000000 452.600000 0.600000 ;
    END
  END psum_norm_1[3]
  PIN psum_norm_1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.600000 0.000000 451.800000 0.600000 ;
    END
  END psum_norm_1[2]
  PIN psum_norm_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.800000 0.000000 451.000000 0.600000 ;
    END
  END psum_norm_1[1]
  PIN psum_norm_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.000000 0.000000 450.200000 0.600000 ;
    END
  END psum_norm_1[0]
  PIN psum_norm_2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.200000 0.000000 449.400000 0.600000 ;
    END
  END psum_norm_2[10]
  PIN psum_norm_2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.400000 0.000000 448.600000 0.600000 ;
    END
  END psum_norm_2[9]
  PIN psum_norm_2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.600000 0.000000 447.800000 0.600000 ;
    END
  END psum_norm_2[8]
  PIN psum_norm_2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.800000 0.000000 447.000000 0.600000 ;
    END
  END psum_norm_2[7]
  PIN psum_norm_2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.000000 0.000000 446.200000 0.600000 ;
    END
  END psum_norm_2[6]
  PIN psum_norm_2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.200000 0.000000 445.400000 0.600000 ;
    END
  END psum_norm_2[5]
  PIN psum_norm_2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.400000 0.000000 444.600000 0.600000 ;
    END
  END psum_norm_2[4]
  PIN psum_norm_2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.600000 0.000000 443.800000 0.600000 ;
    END
  END psum_norm_2[3]
  PIN psum_norm_2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.800000 0.000000 443.000000 0.600000 ;
    END
  END psum_norm_2[2]
  PIN psum_norm_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.000000 0.000000 442.200000 0.600000 ;
    END
  END psum_norm_2[1]
  PIN psum_norm_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.200000 0.000000 441.400000 0.600000 ;
    END
  END psum_norm_2[0]
  PIN norm_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 458.800000 0.000000 459.000000 0.600000 ;
    END
  END norm_valid
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 568.000000 565.400000 ;
    LAYER M2 ;
      RECT 0.000000 0.700000 568.000000 565.400000 ;
      RECT 460.700000 0.000000 568.000000 0.700000 ;
      RECT 459.900000 0.000000 460.300000 0.700000 ;
      RECT 459.100000 0.000000 459.500000 0.700000 ;
      RECT 458.300000 0.000000 458.700000 0.700000 ;
      RECT 457.500000 0.000000 457.900000 0.700000 ;
      RECT 456.700000 0.000000 457.100000 0.700000 ;
      RECT 455.900000 0.000000 456.300000 0.700000 ;
      RECT 455.100000 0.000000 455.500000 0.700000 ;
      RECT 454.300000 0.000000 454.700000 0.700000 ;
      RECT 453.500000 0.000000 453.900000 0.700000 ;
      RECT 452.700000 0.000000 453.100000 0.700000 ;
      RECT 451.900000 0.000000 452.300000 0.700000 ;
      RECT 451.100000 0.000000 451.500000 0.700000 ;
      RECT 450.300000 0.000000 450.700000 0.700000 ;
      RECT 449.500000 0.000000 449.900000 0.700000 ;
      RECT 448.700000 0.000000 449.100000 0.700000 ;
      RECT 447.900000 0.000000 448.300000 0.700000 ;
      RECT 447.100000 0.000000 447.500000 0.700000 ;
      RECT 446.300000 0.000000 446.700000 0.700000 ;
      RECT 445.500000 0.000000 445.900000 0.700000 ;
      RECT 444.700000 0.000000 445.100000 0.700000 ;
      RECT 443.900000 0.000000 444.300000 0.700000 ;
      RECT 443.100000 0.000000 443.500000 0.700000 ;
      RECT 442.300000 0.000000 442.700000 0.700000 ;
      RECT 441.500000 0.000000 441.900000 0.700000 ;
      RECT 440.700000 0.000000 441.100000 0.700000 ;
      RECT 439.900000 0.000000 440.300000 0.700000 ;
      RECT 439.100000 0.000000 439.500000 0.700000 ;
      RECT 438.300000 0.000000 438.700000 0.700000 ;
      RECT 437.500000 0.000000 437.900000 0.700000 ;
      RECT 436.700000 0.000000 437.100000 0.700000 ;
      RECT 435.900000 0.000000 436.300000 0.700000 ;
      RECT 435.100000 0.000000 435.500000 0.700000 ;
      RECT 434.300000 0.000000 434.700000 0.700000 ;
      RECT 433.500000 0.000000 433.900000 0.700000 ;
      RECT 432.700000 0.000000 433.100000 0.700000 ;
      RECT 431.900000 0.000000 432.300000 0.700000 ;
      RECT 431.100000 0.000000 431.500000 0.700000 ;
      RECT 430.300000 0.000000 430.700000 0.700000 ;
      RECT 429.500000 0.000000 429.900000 0.700000 ;
      RECT 428.700000 0.000000 429.100000 0.700000 ;
      RECT 427.900000 0.000000 428.300000 0.700000 ;
      RECT 427.100000 0.000000 427.500000 0.700000 ;
      RECT 426.300000 0.000000 426.700000 0.700000 ;
      RECT 425.500000 0.000000 425.900000 0.700000 ;
      RECT 424.700000 0.000000 425.100000 0.700000 ;
      RECT 423.900000 0.000000 424.300000 0.700000 ;
      RECT 423.100000 0.000000 423.500000 0.700000 ;
      RECT 422.300000 0.000000 422.700000 0.700000 ;
      RECT 421.500000 0.000000 421.900000 0.700000 ;
      RECT 420.700000 0.000000 421.100000 0.700000 ;
      RECT 419.900000 0.000000 420.300000 0.700000 ;
      RECT 419.100000 0.000000 419.500000 0.700000 ;
      RECT 418.300000 0.000000 418.700000 0.700000 ;
      RECT 417.500000 0.000000 417.900000 0.700000 ;
      RECT 416.700000 0.000000 417.100000 0.700000 ;
      RECT 415.900000 0.000000 416.300000 0.700000 ;
      RECT 415.100000 0.000000 415.500000 0.700000 ;
      RECT 414.300000 0.000000 414.700000 0.700000 ;
      RECT 413.500000 0.000000 413.900000 0.700000 ;
      RECT 412.700000 0.000000 413.100000 0.700000 ;
      RECT 411.900000 0.000000 412.300000 0.700000 ;
      RECT 411.100000 0.000000 411.500000 0.700000 ;
      RECT 410.300000 0.000000 410.700000 0.700000 ;
      RECT 409.500000 0.000000 409.900000 0.700000 ;
      RECT 408.700000 0.000000 409.100000 0.700000 ;
      RECT 407.900000 0.000000 408.300000 0.700000 ;
      RECT 407.100000 0.000000 407.500000 0.700000 ;
      RECT 406.300000 0.000000 406.700000 0.700000 ;
      RECT 405.500000 0.000000 405.900000 0.700000 ;
      RECT 404.700000 0.000000 405.100000 0.700000 ;
      RECT 403.900000 0.000000 404.300000 0.700000 ;
      RECT 403.100000 0.000000 403.500000 0.700000 ;
      RECT 402.300000 0.000000 402.700000 0.700000 ;
      RECT 401.500000 0.000000 401.900000 0.700000 ;
      RECT 400.700000 0.000000 401.100000 0.700000 ;
      RECT 399.900000 0.000000 400.300000 0.700000 ;
      RECT 399.100000 0.000000 399.500000 0.700000 ;
      RECT 398.300000 0.000000 398.700000 0.700000 ;
      RECT 397.500000 0.000000 397.900000 0.700000 ;
      RECT 396.700000 0.000000 397.100000 0.700000 ;
      RECT 395.900000 0.000000 396.300000 0.700000 ;
      RECT 395.100000 0.000000 395.500000 0.700000 ;
      RECT 394.300000 0.000000 394.700000 0.700000 ;
      RECT 393.500000 0.000000 393.900000 0.700000 ;
      RECT 392.700000 0.000000 393.100000 0.700000 ;
      RECT 391.900000 0.000000 392.300000 0.700000 ;
      RECT 391.100000 0.000000 391.500000 0.700000 ;
      RECT 390.300000 0.000000 390.700000 0.700000 ;
      RECT 389.500000 0.000000 389.900000 0.700000 ;
      RECT 388.700000 0.000000 389.100000 0.700000 ;
      RECT 387.900000 0.000000 388.300000 0.700000 ;
      RECT 387.100000 0.000000 387.500000 0.700000 ;
      RECT 386.300000 0.000000 386.700000 0.700000 ;
      RECT 385.500000 0.000000 385.900000 0.700000 ;
      RECT 384.700000 0.000000 385.100000 0.700000 ;
      RECT 383.900000 0.000000 384.300000 0.700000 ;
      RECT 383.100000 0.000000 383.500000 0.700000 ;
      RECT 382.300000 0.000000 382.700000 0.700000 ;
      RECT 381.500000 0.000000 381.900000 0.700000 ;
      RECT 380.700000 0.000000 381.100000 0.700000 ;
      RECT 379.900000 0.000000 380.300000 0.700000 ;
      RECT 379.100000 0.000000 379.500000 0.700000 ;
      RECT 378.300000 0.000000 378.700000 0.700000 ;
      RECT 377.500000 0.000000 377.900000 0.700000 ;
      RECT 376.700000 0.000000 377.100000 0.700000 ;
      RECT 375.900000 0.000000 376.300000 0.700000 ;
      RECT 375.100000 0.000000 375.500000 0.700000 ;
      RECT 374.300000 0.000000 374.700000 0.700000 ;
      RECT 373.500000 0.000000 373.900000 0.700000 ;
      RECT 372.700000 0.000000 373.100000 0.700000 ;
      RECT 371.900000 0.000000 372.300000 0.700000 ;
      RECT 371.100000 0.000000 371.500000 0.700000 ;
      RECT 370.300000 0.000000 370.700000 0.700000 ;
      RECT 369.500000 0.000000 369.900000 0.700000 ;
      RECT 368.700000 0.000000 369.100000 0.700000 ;
      RECT 367.900000 0.000000 368.300000 0.700000 ;
      RECT 367.100000 0.000000 367.500000 0.700000 ;
      RECT 366.300000 0.000000 366.700000 0.700000 ;
      RECT 365.500000 0.000000 365.900000 0.700000 ;
      RECT 364.700000 0.000000 365.100000 0.700000 ;
      RECT 363.900000 0.000000 364.300000 0.700000 ;
      RECT 363.100000 0.000000 363.500000 0.700000 ;
      RECT 362.300000 0.000000 362.700000 0.700000 ;
      RECT 361.500000 0.000000 361.900000 0.700000 ;
      RECT 360.700000 0.000000 361.100000 0.700000 ;
      RECT 359.900000 0.000000 360.300000 0.700000 ;
      RECT 359.100000 0.000000 359.500000 0.700000 ;
      RECT 358.300000 0.000000 358.700000 0.700000 ;
      RECT 357.500000 0.000000 357.900000 0.700000 ;
      RECT 356.700000 0.000000 357.100000 0.700000 ;
      RECT 355.900000 0.000000 356.300000 0.700000 ;
      RECT 355.100000 0.000000 355.500000 0.700000 ;
      RECT 354.300000 0.000000 354.700000 0.700000 ;
      RECT 353.500000 0.000000 353.900000 0.700000 ;
      RECT 352.700000 0.000000 353.100000 0.700000 ;
      RECT 351.900000 0.000000 352.300000 0.700000 ;
      RECT 351.100000 0.000000 351.500000 0.700000 ;
      RECT 350.300000 0.000000 350.700000 0.700000 ;
      RECT 349.500000 0.000000 349.900000 0.700000 ;
      RECT 348.700000 0.000000 349.100000 0.700000 ;
      RECT 347.900000 0.000000 348.300000 0.700000 ;
      RECT 347.100000 0.000000 347.500000 0.700000 ;
      RECT 346.300000 0.000000 346.700000 0.700000 ;
      RECT 345.500000 0.000000 345.900000 0.700000 ;
      RECT 344.700000 0.000000 345.100000 0.700000 ;
      RECT 343.900000 0.000000 344.300000 0.700000 ;
      RECT 343.100000 0.000000 343.500000 0.700000 ;
      RECT 342.300000 0.000000 342.700000 0.700000 ;
      RECT 341.500000 0.000000 341.900000 0.700000 ;
      RECT 340.700000 0.000000 341.100000 0.700000 ;
      RECT 339.900000 0.000000 340.300000 0.700000 ;
      RECT 339.100000 0.000000 339.500000 0.700000 ;
      RECT 338.300000 0.000000 338.700000 0.700000 ;
      RECT 337.500000 0.000000 337.900000 0.700000 ;
      RECT 336.700000 0.000000 337.100000 0.700000 ;
      RECT 335.900000 0.000000 336.300000 0.700000 ;
      RECT 335.100000 0.000000 335.500000 0.700000 ;
      RECT 334.300000 0.000000 334.700000 0.700000 ;
      RECT 333.500000 0.000000 333.900000 0.700000 ;
      RECT 332.700000 0.000000 333.100000 0.700000 ;
      RECT 331.900000 0.000000 332.300000 0.700000 ;
      RECT 331.100000 0.000000 331.500000 0.700000 ;
      RECT 330.300000 0.000000 330.700000 0.700000 ;
      RECT 329.500000 0.000000 329.900000 0.700000 ;
      RECT 328.700000 0.000000 329.100000 0.700000 ;
      RECT 327.900000 0.000000 328.300000 0.700000 ;
      RECT 327.100000 0.000000 327.500000 0.700000 ;
      RECT 326.300000 0.000000 326.700000 0.700000 ;
      RECT 325.500000 0.000000 325.900000 0.700000 ;
      RECT 324.700000 0.000000 325.100000 0.700000 ;
      RECT 323.900000 0.000000 324.300000 0.700000 ;
      RECT 323.100000 0.000000 323.500000 0.700000 ;
      RECT 322.300000 0.000000 322.700000 0.700000 ;
      RECT 321.500000 0.000000 321.900000 0.700000 ;
      RECT 320.700000 0.000000 321.100000 0.700000 ;
      RECT 319.900000 0.000000 320.300000 0.700000 ;
      RECT 319.100000 0.000000 319.500000 0.700000 ;
      RECT 318.300000 0.000000 318.700000 0.700000 ;
      RECT 317.500000 0.000000 317.900000 0.700000 ;
      RECT 316.700000 0.000000 317.100000 0.700000 ;
      RECT 315.900000 0.000000 316.300000 0.700000 ;
      RECT 315.100000 0.000000 315.500000 0.700000 ;
      RECT 314.300000 0.000000 314.700000 0.700000 ;
      RECT 313.500000 0.000000 313.900000 0.700000 ;
      RECT 312.700000 0.000000 313.100000 0.700000 ;
      RECT 311.900000 0.000000 312.300000 0.700000 ;
      RECT 311.100000 0.000000 311.500000 0.700000 ;
      RECT 310.300000 0.000000 310.700000 0.700000 ;
      RECT 309.500000 0.000000 309.900000 0.700000 ;
      RECT 308.700000 0.000000 309.100000 0.700000 ;
      RECT 307.900000 0.000000 308.300000 0.700000 ;
      RECT 307.100000 0.000000 307.500000 0.700000 ;
      RECT 306.300000 0.000000 306.700000 0.700000 ;
      RECT 305.500000 0.000000 305.900000 0.700000 ;
      RECT 304.700000 0.000000 305.100000 0.700000 ;
      RECT 303.900000 0.000000 304.300000 0.700000 ;
      RECT 303.100000 0.000000 303.500000 0.700000 ;
      RECT 302.300000 0.000000 302.700000 0.700000 ;
      RECT 301.500000 0.000000 301.900000 0.700000 ;
      RECT 300.700000 0.000000 301.100000 0.700000 ;
      RECT 0.000000 0.000000 300.300000 0.700000 ;
    LAYER M3 ;
      RECT 0.000000 460.800000 568.000000 565.400000 ;
      RECT 0.700000 460.400000 568.000000 460.800000 ;
      RECT 0.000000 460.000000 568.000000 460.400000 ;
      RECT 0.700000 459.600000 568.000000 460.000000 ;
      RECT 0.000000 459.200000 568.000000 459.600000 ;
      RECT 0.700000 458.800000 568.000000 459.200000 ;
      RECT 0.000000 458.400000 568.000000 458.800000 ;
      RECT 0.700000 458.000000 568.000000 458.400000 ;
      RECT 0.000000 457.600000 568.000000 458.000000 ;
      RECT 0.700000 457.200000 568.000000 457.600000 ;
      RECT 0.000000 456.800000 568.000000 457.200000 ;
      RECT 0.700000 456.400000 568.000000 456.800000 ;
      RECT 0.000000 456.000000 568.000000 456.400000 ;
      RECT 0.700000 455.600000 568.000000 456.000000 ;
      RECT 0.000000 455.200000 568.000000 455.600000 ;
      RECT 0.700000 454.800000 568.000000 455.200000 ;
      RECT 0.000000 454.400000 568.000000 454.800000 ;
      RECT 0.700000 454.000000 568.000000 454.400000 ;
      RECT 0.000000 453.600000 568.000000 454.000000 ;
      RECT 0.700000 453.200000 568.000000 453.600000 ;
      RECT 0.000000 452.800000 568.000000 453.200000 ;
      RECT 0.700000 452.400000 568.000000 452.800000 ;
      RECT 0.000000 452.000000 568.000000 452.400000 ;
      RECT 0.700000 451.600000 568.000000 452.000000 ;
      RECT 0.000000 451.200000 568.000000 451.600000 ;
      RECT 0.700000 450.800000 568.000000 451.200000 ;
      RECT 0.000000 450.400000 568.000000 450.800000 ;
      RECT 0.700000 450.000000 568.000000 450.400000 ;
      RECT 0.000000 449.600000 568.000000 450.000000 ;
      RECT 0.700000 449.200000 568.000000 449.600000 ;
      RECT 0.000000 448.800000 568.000000 449.200000 ;
      RECT 0.700000 448.400000 568.000000 448.800000 ;
      RECT 0.000000 448.000000 568.000000 448.400000 ;
      RECT 0.700000 447.600000 568.000000 448.000000 ;
      RECT 0.000000 447.200000 568.000000 447.600000 ;
      RECT 0.700000 446.800000 568.000000 447.200000 ;
      RECT 0.000000 446.400000 568.000000 446.800000 ;
      RECT 0.700000 446.000000 568.000000 446.400000 ;
      RECT 0.000000 445.600000 568.000000 446.000000 ;
      RECT 0.700000 445.200000 568.000000 445.600000 ;
      RECT 0.000000 444.800000 568.000000 445.200000 ;
      RECT 0.700000 444.400000 568.000000 444.800000 ;
      RECT 0.000000 444.000000 568.000000 444.400000 ;
      RECT 0.700000 443.600000 568.000000 444.000000 ;
      RECT 0.000000 443.200000 568.000000 443.600000 ;
      RECT 0.700000 442.800000 568.000000 443.200000 ;
      RECT 0.000000 442.400000 568.000000 442.800000 ;
      RECT 0.700000 442.000000 568.000000 442.400000 ;
      RECT 0.000000 441.600000 568.000000 442.000000 ;
      RECT 0.700000 441.200000 568.000000 441.600000 ;
      RECT 0.000000 440.800000 568.000000 441.200000 ;
      RECT 0.700000 440.400000 568.000000 440.800000 ;
      RECT 0.000000 440.000000 568.000000 440.400000 ;
      RECT 0.700000 439.600000 568.000000 440.000000 ;
      RECT 0.000000 439.200000 568.000000 439.600000 ;
      RECT 0.700000 438.800000 568.000000 439.200000 ;
      RECT 0.000000 438.400000 568.000000 438.800000 ;
      RECT 0.700000 438.000000 568.000000 438.400000 ;
      RECT 0.000000 437.600000 568.000000 438.000000 ;
      RECT 0.700000 437.200000 568.000000 437.600000 ;
      RECT 0.000000 436.800000 568.000000 437.200000 ;
      RECT 0.700000 436.400000 568.000000 436.800000 ;
      RECT 0.000000 436.000000 568.000000 436.400000 ;
      RECT 0.700000 435.600000 568.000000 436.000000 ;
      RECT 0.000000 435.200000 568.000000 435.600000 ;
      RECT 0.700000 434.800000 568.000000 435.200000 ;
      RECT 0.000000 434.400000 568.000000 434.800000 ;
      RECT 0.700000 434.000000 568.000000 434.400000 ;
      RECT 0.000000 433.600000 568.000000 434.000000 ;
      RECT 0.700000 433.200000 568.000000 433.600000 ;
      RECT 0.000000 432.800000 568.000000 433.200000 ;
      RECT 0.700000 432.400000 568.000000 432.800000 ;
      RECT 0.000000 432.000000 568.000000 432.400000 ;
      RECT 0.700000 431.600000 568.000000 432.000000 ;
      RECT 0.000000 431.200000 568.000000 431.600000 ;
      RECT 0.700000 430.800000 568.000000 431.200000 ;
      RECT 0.000000 430.400000 568.000000 430.800000 ;
      RECT 0.700000 430.000000 568.000000 430.400000 ;
      RECT 0.000000 429.600000 568.000000 430.000000 ;
      RECT 0.700000 429.200000 568.000000 429.600000 ;
      RECT 0.000000 428.800000 568.000000 429.200000 ;
      RECT 0.700000 428.400000 568.000000 428.800000 ;
      RECT 0.000000 428.000000 568.000000 428.400000 ;
      RECT 0.700000 427.600000 568.000000 428.000000 ;
      RECT 0.000000 427.200000 568.000000 427.600000 ;
      RECT 0.700000 426.800000 568.000000 427.200000 ;
      RECT 0.000000 426.400000 568.000000 426.800000 ;
      RECT 0.700000 426.000000 568.000000 426.400000 ;
      RECT 0.000000 425.600000 568.000000 426.000000 ;
      RECT 0.700000 425.200000 568.000000 425.600000 ;
      RECT 0.000000 424.800000 568.000000 425.200000 ;
      RECT 0.700000 424.400000 568.000000 424.800000 ;
      RECT 0.000000 424.000000 568.000000 424.400000 ;
      RECT 0.700000 423.600000 568.000000 424.000000 ;
      RECT 0.000000 423.200000 568.000000 423.600000 ;
      RECT 0.700000 422.800000 568.000000 423.200000 ;
      RECT 0.000000 422.400000 568.000000 422.800000 ;
      RECT 0.700000 422.000000 568.000000 422.400000 ;
      RECT 0.000000 421.600000 568.000000 422.000000 ;
      RECT 0.700000 421.200000 568.000000 421.600000 ;
      RECT 0.000000 420.800000 568.000000 421.200000 ;
      RECT 0.700000 420.400000 568.000000 420.800000 ;
      RECT 0.000000 420.000000 568.000000 420.400000 ;
      RECT 0.700000 419.600000 568.000000 420.000000 ;
      RECT 0.000000 419.200000 568.000000 419.600000 ;
      RECT 0.700000 418.800000 568.000000 419.200000 ;
      RECT 0.000000 418.400000 568.000000 418.800000 ;
      RECT 0.700000 418.000000 568.000000 418.400000 ;
      RECT 0.000000 417.600000 568.000000 418.000000 ;
      RECT 0.700000 417.200000 568.000000 417.600000 ;
      RECT 0.000000 416.800000 568.000000 417.200000 ;
      RECT 0.700000 416.400000 568.000000 416.800000 ;
      RECT 0.000000 416.000000 568.000000 416.400000 ;
      RECT 0.700000 415.600000 568.000000 416.000000 ;
      RECT 0.000000 415.200000 568.000000 415.600000 ;
      RECT 0.700000 414.800000 568.000000 415.200000 ;
      RECT 0.000000 414.400000 568.000000 414.800000 ;
      RECT 0.700000 414.000000 568.000000 414.400000 ;
      RECT 0.000000 413.600000 568.000000 414.000000 ;
      RECT 0.700000 413.200000 568.000000 413.600000 ;
      RECT 0.000000 412.800000 568.000000 413.200000 ;
      RECT 0.700000 412.400000 568.000000 412.800000 ;
      RECT 0.000000 412.000000 568.000000 412.400000 ;
      RECT 0.700000 411.600000 568.000000 412.000000 ;
      RECT 0.000000 411.200000 568.000000 411.600000 ;
      RECT 0.700000 410.800000 568.000000 411.200000 ;
      RECT 0.000000 410.400000 568.000000 410.800000 ;
      RECT 0.700000 410.000000 568.000000 410.400000 ;
      RECT 0.000000 409.600000 568.000000 410.000000 ;
      RECT 0.700000 409.200000 568.000000 409.600000 ;
      RECT 0.000000 408.800000 568.000000 409.200000 ;
      RECT 0.700000 408.400000 568.000000 408.800000 ;
      RECT 0.000000 408.000000 568.000000 408.400000 ;
      RECT 0.700000 407.600000 568.000000 408.000000 ;
      RECT 0.000000 407.200000 568.000000 407.600000 ;
      RECT 0.700000 406.800000 568.000000 407.200000 ;
      RECT 0.000000 406.400000 568.000000 406.800000 ;
      RECT 0.700000 406.000000 568.000000 406.400000 ;
      RECT 0.000000 405.600000 568.000000 406.000000 ;
      RECT 0.700000 405.200000 568.000000 405.600000 ;
      RECT 0.000000 404.800000 568.000000 405.200000 ;
      RECT 0.700000 404.400000 568.000000 404.800000 ;
      RECT 0.000000 404.000000 568.000000 404.400000 ;
      RECT 0.700000 403.600000 568.000000 404.000000 ;
      RECT 0.000000 403.200000 568.000000 403.600000 ;
      RECT 0.700000 402.800000 568.000000 403.200000 ;
      RECT 0.000000 402.400000 568.000000 402.800000 ;
      RECT 0.700000 402.000000 568.000000 402.400000 ;
      RECT 0.000000 401.600000 568.000000 402.000000 ;
      RECT 0.700000 401.200000 568.000000 401.600000 ;
      RECT 0.000000 400.800000 568.000000 401.200000 ;
      RECT 0.700000 400.400000 568.000000 400.800000 ;
      RECT 0.000000 400.000000 568.000000 400.400000 ;
      RECT 0.700000 399.600000 568.000000 400.000000 ;
      RECT 0.000000 399.200000 568.000000 399.600000 ;
      RECT 0.700000 398.800000 568.000000 399.200000 ;
      RECT 0.000000 398.400000 568.000000 398.800000 ;
      RECT 0.700000 398.000000 568.000000 398.400000 ;
      RECT 0.000000 397.600000 568.000000 398.000000 ;
      RECT 0.700000 397.200000 568.000000 397.600000 ;
      RECT 0.000000 396.800000 568.000000 397.200000 ;
      RECT 0.700000 396.400000 568.000000 396.800000 ;
      RECT 0.000000 396.000000 568.000000 396.400000 ;
      RECT 0.700000 395.600000 568.000000 396.000000 ;
      RECT 0.000000 395.200000 568.000000 395.600000 ;
      RECT 0.700000 394.800000 568.000000 395.200000 ;
      RECT 0.000000 394.400000 568.000000 394.800000 ;
      RECT 0.700000 394.000000 568.000000 394.400000 ;
      RECT 0.000000 393.600000 568.000000 394.000000 ;
      RECT 0.700000 393.200000 568.000000 393.600000 ;
      RECT 0.000000 392.800000 568.000000 393.200000 ;
      RECT 0.700000 392.400000 568.000000 392.800000 ;
      RECT 0.000000 392.000000 568.000000 392.400000 ;
      RECT 0.700000 391.600000 568.000000 392.000000 ;
      RECT 0.000000 391.200000 568.000000 391.600000 ;
      RECT 0.700000 390.800000 568.000000 391.200000 ;
      RECT 0.000000 390.400000 568.000000 390.800000 ;
      RECT 0.700000 390.000000 568.000000 390.400000 ;
      RECT 0.000000 389.600000 568.000000 390.000000 ;
      RECT 0.700000 389.200000 568.000000 389.600000 ;
      RECT 0.000000 388.800000 568.000000 389.200000 ;
      RECT 0.700000 388.400000 568.000000 388.800000 ;
      RECT 0.000000 388.000000 568.000000 388.400000 ;
      RECT 0.700000 387.600000 568.000000 388.000000 ;
      RECT 0.000000 387.200000 568.000000 387.600000 ;
      RECT 0.700000 386.800000 568.000000 387.200000 ;
      RECT 0.000000 386.400000 568.000000 386.800000 ;
      RECT 0.700000 386.000000 568.000000 386.400000 ;
      RECT 0.000000 385.600000 568.000000 386.000000 ;
      RECT 0.700000 385.200000 568.000000 385.600000 ;
      RECT 0.000000 384.800000 568.000000 385.200000 ;
      RECT 0.700000 384.400000 568.000000 384.800000 ;
      RECT 0.000000 384.000000 568.000000 384.400000 ;
      RECT 0.700000 383.600000 568.000000 384.000000 ;
      RECT 0.000000 383.200000 568.000000 383.600000 ;
      RECT 0.700000 382.800000 568.000000 383.200000 ;
      RECT 0.000000 382.400000 568.000000 382.800000 ;
      RECT 0.700000 382.000000 568.000000 382.400000 ;
      RECT 0.000000 381.600000 568.000000 382.000000 ;
      RECT 0.700000 381.200000 568.000000 381.600000 ;
      RECT 0.000000 380.800000 568.000000 381.200000 ;
      RECT 0.700000 380.400000 568.000000 380.800000 ;
      RECT 0.000000 380.000000 568.000000 380.400000 ;
      RECT 0.700000 379.600000 568.000000 380.000000 ;
      RECT 0.000000 379.200000 568.000000 379.600000 ;
      RECT 0.700000 378.800000 568.000000 379.200000 ;
      RECT 0.000000 378.400000 568.000000 378.800000 ;
      RECT 0.700000 378.000000 568.000000 378.400000 ;
      RECT 0.000000 0.000000 568.000000 378.000000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 568.000000 565.400000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 568.000000 565.400000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 568.000000 565.400000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 568.000000 565.400000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 568.000000 565.400000 ;
  END
END dualcore

END LIBRARY
