##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Tue Mar 21 16:03:51 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 441.600000 BY 441.200000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 196.750000 0.600000 196.850000 ;
    END
  END clk
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 243.150000 0.600000 243.250000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 242.350000 0.600000 242.450000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 241.550000 0.600000 241.650000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 240.750000 0.600000 240.850000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 239.950000 0.600000 240.050000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 239.150000 0.600000 239.250000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 238.350000 0.600000 238.450000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 237.550000 0.600000 237.650000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 236.750000 0.600000 236.850000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 235.950000 0.600000 236.050000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 235.150000 0.600000 235.250000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 234.350000 0.600000 234.450000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 233.550000 0.600000 233.650000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 232.750000 0.600000 232.850000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 231.950000 0.600000 232.050000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 231.150000 0.600000 231.250000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 230.350000 0.600000 230.450000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 229.550000 0.600000 229.650000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 228.750000 0.600000 228.850000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 227.950000 0.600000 228.050000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 227.150000 0.600000 227.250000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 226.350000 0.600000 226.450000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 225.550000 0.600000 225.650000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 224.750000 0.600000 224.850000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 223.950000 0.600000 224.050000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 223.150000 0.600000 223.250000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 222.350000 0.600000 222.450000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 221.550000 0.600000 221.650000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 220.750000 0.600000 220.850000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 219.950000 0.600000 220.050000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 219.150000 0.600000 219.250000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 218.350000 0.600000 218.450000 ;
    END
  END mem_in[0]
  PIN inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 217.550000 0.600000 217.650000 ;
    END
  END inst[25]
  PIN inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 216.750000 0.600000 216.850000 ;
    END
  END inst[24]
  PIN inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 215.950000 0.600000 216.050000 ;
    END
  END inst[23]
  PIN inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 215.150000 0.600000 215.250000 ;
    END
  END inst[22]
  PIN inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 214.350000 0.600000 214.450000 ;
    END
  END inst[21]
  PIN inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 213.550000 0.600000 213.650000 ;
    END
  END inst[20]
  PIN inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 212.750000 0.600000 212.850000 ;
    END
  END inst[19]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 211.950000 0.600000 212.050000 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 211.150000 0.600000 211.250000 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 210.350000 0.600000 210.450000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 209.550000 0.600000 209.650000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 208.750000 0.600000 208.850000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 207.950000 0.600000 208.050000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 207.150000 0.600000 207.250000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 206.350000 0.600000 206.450000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 205.550000 0.600000 205.650000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 204.750000 0.600000 204.850000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 203.950000 0.600000 204.050000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 203.150000 0.600000 203.250000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 202.350000 0.600000 202.450000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 201.550000 0.600000 201.650000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 200.750000 0.600000 200.850000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 199.950000 0.600000 200.050000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 199.150000 0.600000 199.250000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 198.350000 0.600000 198.450000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 197.550000 0.600000 197.650000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 243.950000 0.600000 244.050000 ;
    END
  END reset
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 185.950000 441.600000 186.050000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 186.750000 441.600000 186.850000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 187.550000 441.600000 187.650000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 188.350000 441.600000 188.450000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 189.150000 441.600000 189.250000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 189.950000 441.600000 190.050000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 190.750000 441.600000 190.850000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 191.550000 441.600000 191.650000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 192.350000 441.600000 192.450000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 193.150000 441.600000 193.250000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 193.950000 441.600000 194.050000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 194.750000 441.600000 194.850000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 195.550000 441.600000 195.650000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 196.350000 441.600000 196.450000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 197.150000 441.600000 197.250000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 197.950000 441.600000 198.050000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 198.750000 441.600000 198.850000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 199.550000 441.600000 199.650000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 200.350000 441.600000 200.450000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 201.150000 441.600000 201.250000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 201.950000 441.600000 202.050000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 202.750000 441.600000 202.850000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 203.550000 441.600000 203.650000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 204.350000 441.600000 204.450000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 205.150000 441.600000 205.250000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 205.950000 441.600000 206.050000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 206.750000 441.600000 206.850000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 207.550000 441.600000 207.650000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 208.350000 441.600000 208.450000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 209.150000 441.600000 209.250000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 209.950000 441.600000 210.050000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 210.750000 441.600000 210.850000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 211.550000 441.600000 211.650000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 212.350000 441.600000 212.450000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 213.150000 441.600000 213.250000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 213.950000 441.600000 214.050000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 214.750000 441.600000 214.850000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 215.550000 441.600000 215.650000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 216.350000 441.600000 216.450000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 217.150000 441.600000 217.250000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 217.950000 441.600000 218.050000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 218.750000 441.600000 218.850000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 219.550000 441.600000 219.650000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 220.350000 441.600000 220.450000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 221.150000 441.600000 221.250000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 221.950000 441.600000 222.050000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 222.750000 441.600000 222.850000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 223.550000 441.600000 223.650000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 224.350000 441.600000 224.450000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 225.150000 441.600000 225.250000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 225.950000 441.600000 226.050000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 226.750000 441.600000 226.850000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 227.550000 441.600000 227.650000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 228.350000 441.600000 228.450000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 229.150000 441.600000 229.250000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 229.950000 441.600000 230.050000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 230.750000 441.600000 230.850000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 231.550000 441.600000 231.650000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 232.350000 441.600000 232.450000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 233.150000 441.600000 233.250000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 233.950000 441.600000 234.050000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 234.750000 441.600000 234.850000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 235.550000 441.600000 235.650000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 236.350000 441.600000 236.450000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 237.150000 441.600000 237.250000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 237.950000 441.600000 238.050000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 238.750000 441.600000 238.850000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 239.550000 441.600000 239.650000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 240.350000 441.600000 240.450000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 241.150000 441.600000 241.250000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 241.950000 441.600000 242.050000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 242.750000 441.600000 242.850000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 243.550000 441.600000 243.650000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 244.350000 441.600000 244.450000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 245.150000 441.600000 245.250000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 245.950000 441.600000 246.050000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 246.750000 441.600000 246.850000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 247.550000 441.600000 247.650000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 248.350000 441.600000 248.450000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 249.150000 441.600000 249.250000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 249.950000 441.600000 250.050000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 250.750000 441.600000 250.850000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 251.550000 441.600000 251.650000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 252.350000 441.600000 252.450000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 253.150000 441.600000 253.250000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 253.950000 441.600000 254.050000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 254.750000 441.600000 254.850000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 441.000000 255.550000 441.600000 255.650000 ;
    END
  END out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 441.600000 441.200000 ;
    LAYER M2 ;
      RECT 0.000000 0.000000 441.600000 441.200000 ;
    LAYER M3 ;
      RECT 0.000000 255.750000 441.600000 441.200000 ;
      RECT 0.000000 255.450000 440.880000 255.750000 ;
      RECT 0.000000 254.950000 441.600000 255.450000 ;
      RECT 0.000000 254.650000 440.880000 254.950000 ;
      RECT 0.000000 254.150000 441.600000 254.650000 ;
      RECT 0.000000 253.850000 440.880000 254.150000 ;
      RECT 0.000000 253.350000 441.600000 253.850000 ;
      RECT 0.000000 253.050000 440.880000 253.350000 ;
      RECT 0.000000 252.550000 441.600000 253.050000 ;
      RECT 0.000000 252.250000 440.880000 252.550000 ;
      RECT 0.000000 251.750000 441.600000 252.250000 ;
      RECT 0.000000 251.450000 440.880000 251.750000 ;
      RECT 0.000000 250.950000 441.600000 251.450000 ;
      RECT 0.000000 250.650000 440.880000 250.950000 ;
      RECT 0.000000 250.150000 441.600000 250.650000 ;
      RECT 0.000000 249.850000 440.880000 250.150000 ;
      RECT 0.000000 249.350000 441.600000 249.850000 ;
      RECT 0.000000 249.050000 440.880000 249.350000 ;
      RECT 0.000000 248.550000 441.600000 249.050000 ;
      RECT 0.000000 248.250000 440.880000 248.550000 ;
      RECT 0.000000 247.750000 441.600000 248.250000 ;
      RECT 0.000000 247.450000 440.880000 247.750000 ;
      RECT 0.000000 246.950000 441.600000 247.450000 ;
      RECT 0.000000 246.650000 440.880000 246.950000 ;
      RECT 0.000000 246.150000 441.600000 246.650000 ;
      RECT 0.000000 245.850000 440.880000 246.150000 ;
      RECT 0.000000 245.350000 441.600000 245.850000 ;
      RECT 0.000000 245.050000 440.880000 245.350000 ;
      RECT 0.000000 244.550000 441.600000 245.050000 ;
      RECT 0.000000 244.250000 440.880000 244.550000 ;
      RECT 0.000000 244.150000 441.600000 244.250000 ;
      RECT 0.720000 243.850000 441.600000 244.150000 ;
      RECT 0.000000 243.750000 441.600000 243.850000 ;
      RECT 0.000000 243.450000 440.880000 243.750000 ;
      RECT 0.000000 243.350000 441.600000 243.450000 ;
      RECT 0.720000 243.050000 441.600000 243.350000 ;
      RECT 0.000000 242.950000 441.600000 243.050000 ;
      RECT 0.000000 242.650000 440.880000 242.950000 ;
      RECT 0.000000 242.550000 441.600000 242.650000 ;
      RECT 0.720000 242.250000 441.600000 242.550000 ;
      RECT 0.000000 242.150000 441.600000 242.250000 ;
      RECT 0.000000 241.850000 440.880000 242.150000 ;
      RECT 0.000000 241.750000 441.600000 241.850000 ;
      RECT 0.720000 241.450000 441.600000 241.750000 ;
      RECT 0.000000 241.350000 441.600000 241.450000 ;
      RECT 0.000000 241.050000 440.880000 241.350000 ;
      RECT 0.000000 240.950000 441.600000 241.050000 ;
      RECT 0.720000 240.650000 441.600000 240.950000 ;
      RECT 0.000000 240.550000 441.600000 240.650000 ;
      RECT 0.000000 240.250000 440.880000 240.550000 ;
      RECT 0.000000 240.150000 441.600000 240.250000 ;
      RECT 0.720000 239.850000 441.600000 240.150000 ;
      RECT 0.000000 239.750000 441.600000 239.850000 ;
      RECT 0.000000 239.450000 440.880000 239.750000 ;
      RECT 0.000000 239.350000 441.600000 239.450000 ;
      RECT 0.720000 239.050000 441.600000 239.350000 ;
      RECT 0.000000 238.950000 441.600000 239.050000 ;
      RECT 0.000000 238.650000 440.880000 238.950000 ;
      RECT 0.000000 238.550000 441.600000 238.650000 ;
      RECT 0.720000 238.250000 441.600000 238.550000 ;
      RECT 0.000000 238.150000 441.600000 238.250000 ;
      RECT 0.000000 237.850000 440.880000 238.150000 ;
      RECT 0.000000 237.750000 441.600000 237.850000 ;
      RECT 0.720000 237.450000 441.600000 237.750000 ;
      RECT 0.000000 237.350000 441.600000 237.450000 ;
      RECT 0.000000 237.050000 440.880000 237.350000 ;
      RECT 0.000000 236.950000 441.600000 237.050000 ;
      RECT 0.720000 236.650000 441.600000 236.950000 ;
      RECT 0.000000 236.550000 441.600000 236.650000 ;
      RECT 0.000000 236.250000 440.880000 236.550000 ;
      RECT 0.000000 236.150000 441.600000 236.250000 ;
      RECT 0.720000 235.850000 441.600000 236.150000 ;
      RECT 0.000000 235.750000 441.600000 235.850000 ;
      RECT 0.000000 235.450000 440.880000 235.750000 ;
      RECT 0.000000 235.350000 441.600000 235.450000 ;
      RECT 0.720000 235.050000 441.600000 235.350000 ;
      RECT 0.000000 234.950000 441.600000 235.050000 ;
      RECT 0.000000 234.650000 440.880000 234.950000 ;
      RECT 0.000000 234.550000 441.600000 234.650000 ;
      RECT 0.720000 234.250000 441.600000 234.550000 ;
      RECT 0.000000 234.150000 441.600000 234.250000 ;
      RECT 0.000000 233.850000 440.880000 234.150000 ;
      RECT 0.000000 233.750000 441.600000 233.850000 ;
      RECT 0.720000 233.450000 441.600000 233.750000 ;
      RECT 0.000000 233.350000 441.600000 233.450000 ;
      RECT 0.000000 233.050000 440.880000 233.350000 ;
      RECT 0.000000 232.950000 441.600000 233.050000 ;
      RECT 0.720000 232.650000 441.600000 232.950000 ;
      RECT 0.000000 232.550000 441.600000 232.650000 ;
      RECT 0.000000 232.250000 440.880000 232.550000 ;
      RECT 0.000000 232.150000 441.600000 232.250000 ;
      RECT 0.720000 231.850000 441.600000 232.150000 ;
      RECT 0.000000 231.750000 441.600000 231.850000 ;
      RECT 0.000000 231.450000 440.880000 231.750000 ;
      RECT 0.000000 231.350000 441.600000 231.450000 ;
      RECT 0.720000 231.050000 441.600000 231.350000 ;
      RECT 0.000000 230.950000 441.600000 231.050000 ;
      RECT 0.000000 230.650000 440.880000 230.950000 ;
      RECT 0.000000 230.550000 441.600000 230.650000 ;
      RECT 0.720000 230.250000 441.600000 230.550000 ;
      RECT 0.000000 230.150000 441.600000 230.250000 ;
      RECT 0.000000 229.850000 440.880000 230.150000 ;
      RECT 0.000000 229.750000 441.600000 229.850000 ;
      RECT 0.720000 229.450000 441.600000 229.750000 ;
      RECT 0.000000 229.350000 441.600000 229.450000 ;
      RECT 0.000000 229.050000 440.880000 229.350000 ;
      RECT 0.000000 228.950000 441.600000 229.050000 ;
      RECT 0.720000 228.650000 441.600000 228.950000 ;
      RECT 0.000000 228.550000 441.600000 228.650000 ;
      RECT 0.000000 228.250000 440.880000 228.550000 ;
      RECT 0.000000 228.150000 441.600000 228.250000 ;
      RECT 0.720000 227.850000 441.600000 228.150000 ;
      RECT 0.000000 227.750000 441.600000 227.850000 ;
      RECT 0.000000 227.450000 440.880000 227.750000 ;
      RECT 0.000000 227.350000 441.600000 227.450000 ;
      RECT 0.720000 227.050000 441.600000 227.350000 ;
      RECT 0.000000 226.950000 441.600000 227.050000 ;
      RECT 0.000000 226.650000 440.880000 226.950000 ;
      RECT 0.000000 226.550000 441.600000 226.650000 ;
      RECT 0.720000 226.250000 441.600000 226.550000 ;
      RECT 0.000000 226.150000 441.600000 226.250000 ;
      RECT 0.000000 225.850000 440.880000 226.150000 ;
      RECT 0.000000 225.750000 441.600000 225.850000 ;
      RECT 0.720000 225.450000 441.600000 225.750000 ;
      RECT 0.000000 225.350000 441.600000 225.450000 ;
      RECT 0.000000 225.050000 440.880000 225.350000 ;
      RECT 0.000000 224.950000 441.600000 225.050000 ;
      RECT 0.720000 224.650000 441.600000 224.950000 ;
      RECT 0.000000 224.550000 441.600000 224.650000 ;
      RECT 0.000000 224.250000 440.880000 224.550000 ;
      RECT 0.000000 224.150000 441.600000 224.250000 ;
      RECT 0.720000 223.850000 441.600000 224.150000 ;
      RECT 0.000000 223.750000 441.600000 223.850000 ;
      RECT 0.000000 223.450000 440.880000 223.750000 ;
      RECT 0.000000 223.350000 441.600000 223.450000 ;
      RECT 0.720000 223.050000 441.600000 223.350000 ;
      RECT 0.000000 222.950000 441.600000 223.050000 ;
      RECT 0.000000 222.650000 440.880000 222.950000 ;
      RECT 0.000000 222.550000 441.600000 222.650000 ;
      RECT 0.720000 222.250000 441.600000 222.550000 ;
      RECT 0.000000 222.150000 441.600000 222.250000 ;
      RECT 0.000000 221.850000 440.880000 222.150000 ;
      RECT 0.000000 221.750000 441.600000 221.850000 ;
      RECT 0.720000 221.450000 441.600000 221.750000 ;
      RECT 0.000000 221.350000 441.600000 221.450000 ;
      RECT 0.000000 221.050000 440.880000 221.350000 ;
      RECT 0.000000 220.950000 441.600000 221.050000 ;
      RECT 0.720000 220.650000 441.600000 220.950000 ;
      RECT 0.000000 220.550000 441.600000 220.650000 ;
      RECT 0.000000 220.250000 440.880000 220.550000 ;
      RECT 0.000000 220.150000 441.600000 220.250000 ;
      RECT 0.720000 219.850000 441.600000 220.150000 ;
      RECT 0.000000 219.750000 441.600000 219.850000 ;
      RECT 0.000000 219.450000 440.880000 219.750000 ;
      RECT 0.000000 219.350000 441.600000 219.450000 ;
      RECT 0.720000 219.050000 441.600000 219.350000 ;
      RECT 0.000000 218.950000 441.600000 219.050000 ;
      RECT 0.000000 218.650000 440.880000 218.950000 ;
      RECT 0.000000 218.550000 441.600000 218.650000 ;
      RECT 0.720000 218.250000 441.600000 218.550000 ;
      RECT 0.000000 218.150000 441.600000 218.250000 ;
      RECT 0.000000 217.850000 440.880000 218.150000 ;
      RECT 0.000000 217.750000 441.600000 217.850000 ;
      RECT 0.720000 217.450000 441.600000 217.750000 ;
      RECT 0.000000 217.350000 441.600000 217.450000 ;
      RECT 0.000000 217.050000 440.880000 217.350000 ;
      RECT 0.000000 216.950000 441.600000 217.050000 ;
      RECT 0.720000 216.650000 441.600000 216.950000 ;
      RECT 0.000000 216.550000 441.600000 216.650000 ;
      RECT 0.000000 216.250000 440.880000 216.550000 ;
      RECT 0.000000 216.150000 441.600000 216.250000 ;
      RECT 0.720000 215.850000 441.600000 216.150000 ;
      RECT 0.000000 215.750000 441.600000 215.850000 ;
      RECT 0.000000 215.450000 440.880000 215.750000 ;
      RECT 0.000000 215.350000 441.600000 215.450000 ;
      RECT 0.720000 215.050000 441.600000 215.350000 ;
      RECT 0.000000 214.950000 441.600000 215.050000 ;
      RECT 0.000000 214.650000 440.880000 214.950000 ;
      RECT 0.000000 214.550000 441.600000 214.650000 ;
      RECT 0.720000 214.250000 441.600000 214.550000 ;
      RECT 0.000000 214.150000 441.600000 214.250000 ;
      RECT 0.000000 213.850000 440.880000 214.150000 ;
      RECT 0.000000 213.750000 441.600000 213.850000 ;
      RECT 0.720000 213.450000 441.600000 213.750000 ;
      RECT 0.000000 213.350000 441.600000 213.450000 ;
      RECT 0.000000 213.050000 440.880000 213.350000 ;
      RECT 0.000000 212.950000 441.600000 213.050000 ;
      RECT 0.720000 212.650000 441.600000 212.950000 ;
      RECT 0.000000 212.550000 441.600000 212.650000 ;
      RECT 0.000000 212.250000 440.880000 212.550000 ;
      RECT 0.000000 212.150000 441.600000 212.250000 ;
      RECT 0.720000 211.850000 441.600000 212.150000 ;
      RECT 0.000000 211.750000 441.600000 211.850000 ;
      RECT 0.000000 211.450000 440.880000 211.750000 ;
      RECT 0.000000 211.350000 441.600000 211.450000 ;
      RECT 0.720000 211.050000 441.600000 211.350000 ;
      RECT 0.000000 210.950000 441.600000 211.050000 ;
      RECT 0.000000 210.650000 440.880000 210.950000 ;
      RECT 0.000000 210.550000 441.600000 210.650000 ;
      RECT 0.720000 210.250000 441.600000 210.550000 ;
      RECT 0.000000 210.150000 441.600000 210.250000 ;
      RECT 0.000000 209.850000 440.880000 210.150000 ;
      RECT 0.000000 209.750000 441.600000 209.850000 ;
      RECT 0.720000 209.450000 441.600000 209.750000 ;
      RECT 0.000000 209.350000 441.600000 209.450000 ;
      RECT 0.000000 209.050000 440.880000 209.350000 ;
      RECT 0.000000 208.950000 441.600000 209.050000 ;
      RECT 0.720000 208.650000 441.600000 208.950000 ;
      RECT 0.000000 208.550000 441.600000 208.650000 ;
      RECT 0.000000 208.250000 440.880000 208.550000 ;
      RECT 0.000000 208.150000 441.600000 208.250000 ;
      RECT 0.720000 207.850000 441.600000 208.150000 ;
      RECT 0.000000 207.750000 441.600000 207.850000 ;
      RECT 0.000000 207.450000 440.880000 207.750000 ;
      RECT 0.000000 207.350000 441.600000 207.450000 ;
      RECT 0.720000 207.050000 441.600000 207.350000 ;
      RECT 0.000000 206.950000 441.600000 207.050000 ;
      RECT 0.000000 206.650000 440.880000 206.950000 ;
      RECT 0.000000 206.550000 441.600000 206.650000 ;
      RECT 0.720000 206.250000 441.600000 206.550000 ;
      RECT 0.000000 206.150000 441.600000 206.250000 ;
      RECT 0.000000 205.850000 440.880000 206.150000 ;
      RECT 0.000000 205.750000 441.600000 205.850000 ;
      RECT 0.720000 205.450000 441.600000 205.750000 ;
      RECT 0.000000 205.350000 441.600000 205.450000 ;
      RECT 0.000000 205.050000 440.880000 205.350000 ;
      RECT 0.000000 204.950000 441.600000 205.050000 ;
      RECT 0.720000 204.650000 441.600000 204.950000 ;
      RECT 0.000000 204.550000 441.600000 204.650000 ;
      RECT 0.000000 204.250000 440.880000 204.550000 ;
      RECT 0.000000 204.150000 441.600000 204.250000 ;
      RECT 0.720000 203.850000 441.600000 204.150000 ;
      RECT 0.000000 203.750000 441.600000 203.850000 ;
      RECT 0.000000 203.450000 440.880000 203.750000 ;
      RECT 0.000000 203.350000 441.600000 203.450000 ;
      RECT 0.720000 203.050000 441.600000 203.350000 ;
      RECT 0.000000 202.950000 441.600000 203.050000 ;
      RECT 0.000000 202.650000 440.880000 202.950000 ;
      RECT 0.000000 202.550000 441.600000 202.650000 ;
      RECT 0.720000 202.250000 441.600000 202.550000 ;
      RECT 0.000000 202.150000 441.600000 202.250000 ;
      RECT 0.000000 201.850000 440.880000 202.150000 ;
      RECT 0.000000 201.750000 441.600000 201.850000 ;
      RECT 0.720000 201.450000 441.600000 201.750000 ;
      RECT 0.000000 201.350000 441.600000 201.450000 ;
      RECT 0.000000 201.050000 440.880000 201.350000 ;
      RECT 0.000000 200.950000 441.600000 201.050000 ;
      RECT 0.720000 200.650000 441.600000 200.950000 ;
      RECT 0.000000 200.550000 441.600000 200.650000 ;
      RECT 0.000000 200.250000 440.880000 200.550000 ;
      RECT 0.000000 200.150000 441.600000 200.250000 ;
      RECT 0.720000 199.850000 441.600000 200.150000 ;
      RECT 0.000000 199.750000 441.600000 199.850000 ;
      RECT 0.000000 199.450000 440.880000 199.750000 ;
      RECT 0.000000 199.350000 441.600000 199.450000 ;
      RECT 0.720000 199.050000 441.600000 199.350000 ;
      RECT 0.000000 198.950000 441.600000 199.050000 ;
      RECT 0.000000 198.650000 440.880000 198.950000 ;
      RECT 0.000000 198.550000 441.600000 198.650000 ;
      RECT 0.720000 198.250000 441.600000 198.550000 ;
      RECT 0.000000 198.150000 441.600000 198.250000 ;
      RECT 0.000000 197.850000 440.880000 198.150000 ;
      RECT 0.000000 197.750000 441.600000 197.850000 ;
      RECT 0.720000 197.450000 441.600000 197.750000 ;
      RECT 0.000000 197.350000 441.600000 197.450000 ;
      RECT 0.000000 197.050000 440.880000 197.350000 ;
      RECT 0.000000 196.950000 441.600000 197.050000 ;
      RECT 0.720000 196.650000 441.600000 196.950000 ;
      RECT 0.000000 196.550000 441.600000 196.650000 ;
      RECT 0.000000 196.250000 440.880000 196.550000 ;
      RECT 0.000000 195.750000 441.600000 196.250000 ;
      RECT 0.000000 195.450000 440.880000 195.750000 ;
      RECT 0.000000 194.950000 441.600000 195.450000 ;
      RECT 0.000000 194.650000 440.880000 194.950000 ;
      RECT 0.000000 194.150000 441.600000 194.650000 ;
      RECT 0.000000 193.850000 440.880000 194.150000 ;
      RECT 0.000000 193.350000 441.600000 193.850000 ;
      RECT 0.000000 193.050000 440.880000 193.350000 ;
      RECT 0.000000 192.550000 441.600000 193.050000 ;
      RECT 0.000000 192.250000 440.880000 192.550000 ;
      RECT 0.000000 191.750000 441.600000 192.250000 ;
      RECT 0.000000 191.450000 440.880000 191.750000 ;
      RECT 0.000000 190.950000 441.600000 191.450000 ;
      RECT 0.000000 190.650000 440.880000 190.950000 ;
      RECT 0.000000 190.150000 441.600000 190.650000 ;
      RECT 0.000000 189.850000 440.880000 190.150000 ;
      RECT 0.000000 189.350000 441.600000 189.850000 ;
      RECT 0.000000 189.050000 440.880000 189.350000 ;
      RECT 0.000000 188.550000 441.600000 189.050000 ;
      RECT 0.000000 188.250000 440.880000 188.550000 ;
      RECT 0.000000 187.750000 441.600000 188.250000 ;
      RECT 0.000000 187.450000 440.880000 187.750000 ;
      RECT 0.000000 186.950000 441.600000 187.450000 ;
      RECT 0.000000 186.650000 440.880000 186.950000 ;
      RECT 0.000000 186.150000 441.600000 186.650000 ;
      RECT 0.000000 185.850000 440.880000 186.150000 ;
      RECT 0.000000 0.000000 441.600000 185.850000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 441.600000 441.200000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 441.600000 441.200000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 441.600000 441.200000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 441.600000 441.200000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 441.600000 441.200000 ;
  END
END fullchip

END LIBRARY
