##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Mon Mar 13 01:33:59 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 383.200000 BY 381.800000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 170.750000 0.600000 170.850000 ;
    END
  END clk
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 209.950000 0.600000 210.050000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 209.150000 0.600000 209.250000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 208.350000 0.600000 208.450000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 207.550000 0.600000 207.650000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 206.750000 0.600000 206.850000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 205.950000 0.600000 206.050000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 205.150000 0.600000 205.250000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 204.350000 0.600000 204.450000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 203.550000 0.600000 203.650000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 202.750000 0.600000 202.850000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 201.950000 0.600000 202.050000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 201.150000 0.600000 201.250000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 200.350000 0.600000 200.450000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 199.550000 0.600000 199.650000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 198.750000 0.600000 198.850000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 197.950000 0.600000 198.050000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 197.150000 0.600000 197.250000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 196.350000 0.600000 196.450000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 195.550000 0.600000 195.650000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 194.750000 0.600000 194.850000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 193.950000 0.600000 194.050000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 193.150000 0.600000 193.250000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 192.350000 0.600000 192.450000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 191.550000 0.600000 191.650000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 190.750000 0.600000 190.850000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 189.950000 0.600000 190.050000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 189.150000 0.600000 189.250000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 188.350000 0.600000 188.450000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 187.550000 0.600000 187.650000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 186.750000 0.600000 186.850000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 185.950000 0.600000 186.050000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 185.150000 0.600000 185.250000 ;
    END
  END mem_in[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 184.350000 0.600000 184.450000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 183.550000 0.600000 183.650000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 182.750000 0.600000 182.850000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 181.950000 0.600000 182.050000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 181.150000 0.600000 181.250000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 180.350000 0.600000 180.450000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 179.550000 0.600000 179.650000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 178.750000 0.600000 178.850000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 177.950000 0.600000 178.050000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 177.150000 0.600000 177.250000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 176.350000 0.600000 176.450000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 175.550000 0.600000 175.650000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 174.750000 0.600000 174.850000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 173.950000 0.600000 174.050000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 173.150000 0.600000 173.250000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 172.350000 0.600000 172.450000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 171.550000 0.600000 171.650000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 210.750000 0.600000 210.850000 ;
    END
  END reset
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 156.150000 383.200000 156.250000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 156.950000 383.200000 157.050000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 157.750000 383.200000 157.850000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 158.550000 383.200000 158.650000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 159.350000 383.200000 159.450000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 160.150000 383.200000 160.250000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 160.950000 383.200000 161.050000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 161.750000 383.200000 161.850000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 162.550000 383.200000 162.650000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 163.350000 383.200000 163.450000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 164.150000 383.200000 164.250000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 164.950000 383.200000 165.050000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 165.750000 383.200000 165.850000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 166.550000 383.200000 166.650000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 167.350000 383.200000 167.450000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 168.150000 383.200000 168.250000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 168.950000 383.200000 169.050000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 169.750000 383.200000 169.850000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 170.550000 383.200000 170.650000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 171.350000 383.200000 171.450000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 172.150000 383.200000 172.250000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 172.950000 383.200000 173.050000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 173.750000 383.200000 173.850000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 174.550000 383.200000 174.650000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 175.350000 383.200000 175.450000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 176.150000 383.200000 176.250000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 176.950000 383.200000 177.050000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 177.750000 383.200000 177.850000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 178.550000 383.200000 178.650000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 179.350000 383.200000 179.450000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 180.150000 383.200000 180.250000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 180.950000 383.200000 181.050000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 181.750000 383.200000 181.850000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 182.550000 383.200000 182.650000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 183.350000 383.200000 183.450000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 184.150000 383.200000 184.250000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 184.950000 383.200000 185.050000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 185.750000 383.200000 185.850000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 186.550000 383.200000 186.650000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 187.350000 383.200000 187.450000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 188.150000 383.200000 188.250000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 188.950000 383.200000 189.050000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 189.750000 383.200000 189.850000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 190.550000 383.200000 190.650000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 191.350000 383.200000 191.450000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 192.150000 383.200000 192.250000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 192.950000 383.200000 193.050000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 193.750000 383.200000 193.850000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 194.550000 383.200000 194.650000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 195.350000 383.200000 195.450000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 196.150000 383.200000 196.250000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 196.950000 383.200000 197.050000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 197.750000 383.200000 197.850000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 198.550000 383.200000 198.650000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 199.350000 383.200000 199.450000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 200.150000 383.200000 200.250000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 200.950000 383.200000 201.050000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 201.750000 383.200000 201.850000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 202.550000 383.200000 202.650000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 203.350000 383.200000 203.450000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 204.150000 383.200000 204.250000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 204.950000 383.200000 205.050000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 205.750000 383.200000 205.850000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 206.550000 383.200000 206.650000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 207.350000 383.200000 207.450000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 208.150000 383.200000 208.250000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 208.950000 383.200000 209.050000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 209.750000 383.200000 209.850000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 210.550000 383.200000 210.650000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 211.350000 383.200000 211.450000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 212.150000 383.200000 212.250000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 212.950000 383.200000 213.050000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 213.750000 383.200000 213.850000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 214.550000 383.200000 214.650000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 215.350000 383.200000 215.450000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 216.150000 383.200000 216.250000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 216.950000 383.200000 217.050000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 217.750000 383.200000 217.850000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 218.550000 383.200000 218.650000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 219.350000 383.200000 219.450000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 220.150000 383.200000 220.250000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 220.950000 383.200000 221.050000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 221.750000 383.200000 221.850000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 222.550000 383.200000 222.650000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 223.350000 383.200000 223.450000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 224.150000 383.200000 224.250000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 224.950000 383.200000 225.050000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.600000 225.750000 383.200000 225.850000 ;
    END
  END out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 383.200000 381.800000 ;
    LAYER M2 ;
      RECT 0.000000 0.000000 383.200000 381.800000 ;
    LAYER M3 ;
      RECT 0.000000 225.950000 383.200000 381.800000 ;
      RECT 0.000000 225.650000 382.480000 225.950000 ;
      RECT 0.000000 225.150000 383.200000 225.650000 ;
      RECT 0.000000 224.850000 382.480000 225.150000 ;
      RECT 0.000000 224.350000 383.200000 224.850000 ;
      RECT 0.000000 224.050000 382.480000 224.350000 ;
      RECT 0.000000 223.550000 383.200000 224.050000 ;
      RECT 0.000000 223.250000 382.480000 223.550000 ;
      RECT 0.000000 222.750000 383.200000 223.250000 ;
      RECT 0.000000 222.450000 382.480000 222.750000 ;
      RECT 0.000000 221.950000 383.200000 222.450000 ;
      RECT 0.000000 221.650000 382.480000 221.950000 ;
      RECT 0.000000 221.150000 383.200000 221.650000 ;
      RECT 0.000000 220.850000 382.480000 221.150000 ;
      RECT 0.000000 220.350000 383.200000 220.850000 ;
      RECT 0.000000 220.050000 382.480000 220.350000 ;
      RECT 0.000000 219.550000 383.200000 220.050000 ;
      RECT 0.000000 219.250000 382.480000 219.550000 ;
      RECT 0.000000 218.750000 383.200000 219.250000 ;
      RECT 0.000000 218.450000 382.480000 218.750000 ;
      RECT 0.000000 217.950000 383.200000 218.450000 ;
      RECT 0.000000 217.650000 382.480000 217.950000 ;
      RECT 0.000000 217.150000 383.200000 217.650000 ;
      RECT 0.000000 216.850000 382.480000 217.150000 ;
      RECT 0.000000 216.350000 383.200000 216.850000 ;
      RECT 0.000000 216.050000 382.480000 216.350000 ;
      RECT 0.000000 215.550000 383.200000 216.050000 ;
      RECT 0.000000 215.250000 382.480000 215.550000 ;
      RECT 0.000000 214.750000 383.200000 215.250000 ;
      RECT 0.000000 214.450000 382.480000 214.750000 ;
      RECT 0.000000 213.950000 383.200000 214.450000 ;
      RECT 0.000000 213.650000 382.480000 213.950000 ;
      RECT 0.000000 213.150000 383.200000 213.650000 ;
      RECT 0.000000 212.850000 382.480000 213.150000 ;
      RECT 0.000000 212.350000 383.200000 212.850000 ;
      RECT 0.000000 212.050000 382.480000 212.350000 ;
      RECT 0.000000 211.550000 383.200000 212.050000 ;
      RECT 0.000000 211.250000 382.480000 211.550000 ;
      RECT 0.000000 210.950000 383.200000 211.250000 ;
      RECT 0.720000 210.750000 383.200000 210.950000 ;
      RECT 0.720000 210.650000 382.480000 210.750000 ;
      RECT 0.000000 210.450000 382.480000 210.650000 ;
      RECT 0.000000 210.150000 383.200000 210.450000 ;
      RECT 0.720000 209.950000 383.200000 210.150000 ;
      RECT 0.720000 209.850000 382.480000 209.950000 ;
      RECT 0.000000 209.650000 382.480000 209.850000 ;
      RECT 0.000000 209.350000 383.200000 209.650000 ;
      RECT 0.720000 209.150000 383.200000 209.350000 ;
      RECT 0.720000 209.050000 382.480000 209.150000 ;
      RECT 0.000000 208.850000 382.480000 209.050000 ;
      RECT 0.000000 208.550000 383.200000 208.850000 ;
      RECT 0.720000 208.350000 383.200000 208.550000 ;
      RECT 0.720000 208.250000 382.480000 208.350000 ;
      RECT 0.000000 208.050000 382.480000 208.250000 ;
      RECT 0.000000 207.750000 383.200000 208.050000 ;
      RECT 0.720000 207.550000 383.200000 207.750000 ;
      RECT 0.720000 207.450000 382.480000 207.550000 ;
      RECT 0.000000 207.250000 382.480000 207.450000 ;
      RECT 0.000000 206.950000 383.200000 207.250000 ;
      RECT 0.720000 206.750000 383.200000 206.950000 ;
      RECT 0.720000 206.650000 382.480000 206.750000 ;
      RECT 0.000000 206.450000 382.480000 206.650000 ;
      RECT 0.000000 206.150000 383.200000 206.450000 ;
      RECT 0.720000 205.950000 383.200000 206.150000 ;
      RECT 0.720000 205.850000 382.480000 205.950000 ;
      RECT 0.000000 205.650000 382.480000 205.850000 ;
      RECT 0.000000 205.350000 383.200000 205.650000 ;
      RECT 0.720000 205.150000 383.200000 205.350000 ;
      RECT 0.720000 205.050000 382.480000 205.150000 ;
      RECT 0.000000 204.850000 382.480000 205.050000 ;
      RECT 0.000000 204.550000 383.200000 204.850000 ;
      RECT 0.720000 204.350000 383.200000 204.550000 ;
      RECT 0.720000 204.250000 382.480000 204.350000 ;
      RECT 0.000000 204.050000 382.480000 204.250000 ;
      RECT 0.000000 203.750000 383.200000 204.050000 ;
      RECT 0.720000 203.550000 383.200000 203.750000 ;
      RECT 0.720000 203.450000 382.480000 203.550000 ;
      RECT 0.000000 203.250000 382.480000 203.450000 ;
      RECT 0.000000 202.950000 383.200000 203.250000 ;
      RECT 0.720000 202.750000 383.200000 202.950000 ;
      RECT 0.720000 202.650000 382.480000 202.750000 ;
      RECT 0.000000 202.450000 382.480000 202.650000 ;
      RECT 0.000000 202.150000 383.200000 202.450000 ;
      RECT 0.720000 201.950000 383.200000 202.150000 ;
      RECT 0.720000 201.850000 382.480000 201.950000 ;
      RECT 0.000000 201.650000 382.480000 201.850000 ;
      RECT 0.000000 201.350000 383.200000 201.650000 ;
      RECT 0.720000 201.150000 383.200000 201.350000 ;
      RECT 0.720000 201.050000 382.480000 201.150000 ;
      RECT 0.000000 200.850000 382.480000 201.050000 ;
      RECT 0.000000 200.550000 383.200000 200.850000 ;
      RECT 0.720000 200.350000 383.200000 200.550000 ;
      RECT 0.720000 200.250000 382.480000 200.350000 ;
      RECT 0.000000 200.050000 382.480000 200.250000 ;
      RECT 0.000000 199.750000 383.200000 200.050000 ;
      RECT 0.720000 199.550000 383.200000 199.750000 ;
      RECT 0.720000 199.450000 382.480000 199.550000 ;
      RECT 0.000000 199.250000 382.480000 199.450000 ;
      RECT 0.000000 198.950000 383.200000 199.250000 ;
      RECT 0.720000 198.750000 383.200000 198.950000 ;
      RECT 0.720000 198.650000 382.480000 198.750000 ;
      RECT 0.000000 198.450000 382.480000 198.650000 ;
      RECT 0.000000 198.150000 383.200000 198.450000 ;
      RECT 0.720000 197.950000 383.200000 198.150000 ;
      RECT 0.720000 197.850000 382.480000 197.950000 ;
      RECT 0.000000 197.650000 382.480000 197.850000 ;
      RECT 0.000000 197.350000 383.200000 197.650000 ;
      RECT 0.720000 197.150000 383.200000 197.350000 ;
      RECT 0.720000 197.050000 382.480000 197.150000 ;
      RECT 0.000000 196.850000 382.480000 197.050000 ;
      RECT 0.000000 196.550000 383.200000 196.850000 ;
      RECT 0.720000 196.350000 383.200000 196.550000 ;
      RECT 0.720000 196.250000 382.480000 196.350000 ;
      RECT 0.000000 196.050000 382.480000 196.250000 ;
      RECT 0.000000 195.750000 383.200000 196.050000 ;
      RECT 0.720000 195.550000 383.200000 195.750000 ;
      RECT 0.720000 195.450000 382.480000 195.550000 ;
      RECT 0.000000 195.250000 382.480000 195.450000 ;
      RECT 0.000000 194.950000 383.200000 195.250000 ;
      RECT 0.720000 194.750000 383.200000 194.950000 ;
      RECT 0.720000 194.650000 382.480000 194.750000 ;
      RECT 0.000000 194.450000 382.480000 194.650000 ;
      RECT 0.000000 194.150000 383.200000 194.450000 ;
      RECT 0.720000 193.950000 383.200000 194.150000 ;
      RECT 0.720000 193.850000 382.480000 193.950000 ;
      RECT 0.000000 193.650000 382.480000 193.850000 ;
      RECT 0.000000 193.350000 383.200000 193.650000 ;
      RECT 0.720000 193.150000 383.200000 193.350000 ;
      RECT 0.720000 193.050000 382.480000 193.150000 ;
      RECT 0.000000 192.850000 382.480000 193.050000 ;
      RECT 0.000000 192.550000 383.200000 192.850000 ;
      RECT 0.720000 192.350000 383.200000 192.550000 ;
      RECT 0.720000 192.250000 382.480000 192.350000 ;
      RECT 0.000000 192.050000 382.480000 192.250000 ;
      RECT 0.000000 191.750000 383.200000 192.050000 ;
      RECT 0.720000 191.550000 383.200000 191.750000 ;
      RECT 0.720000 191.450000 382.480000 191.550000 ;
      RECT 0.000000 191.250000 382.480000 191.450000 ;
      RECT 0.000000 190.950000 383.200000 191.250000 ;
      RECT 0.720000 190.750000 383.200000 190.950000 ;
      RECT 0.720000 190.650000 382.480000 190.750000 ;
      RECT 0.000000 190.450000 382.480000 190.650000 ;
      RECT 0.000000 190.150000 383.200000 190.450000 ;
      RECT 0.720000 189.950000 383.200000 190.150000 ;
      RECT 0.720000 189.850000 382.480000 189.950000 ;
      RECT 0.000000 189.650000 382.480000 189.850000 ;
      RECT 0.000000 189.350000 383.200000 189.650000 ;
      RECT 0.720000 189.150000 383.200000 189.350000 ;
      RECT 0.720000 189.050000 382.480000 189.150000 ;
      RECT 0.000000 188.850000 382.480000 189.050000 ;
      RECT 0.000000 188.550000 383.200000 188.850000 ;
      RECT 0.720000 188.350000 383.200000 188.550000 ;
      RECT 0.720000 188.250000 382.480000 188.350000 ;
      RECT 0.000000 188.050000 382.480000 188.250000 ;
      RECT 0.000000 187.750000 383.200000 188.050000 ;
      RECT 0.720000 187.550000 383.200000 187.750000 ;
      RECT 0.720000 187.450000 382.480000 187.550000 ;
      RECT 0.000000 187.250000 382.480000 187.450000 ;
      RECT 0.000000 186.950000 383.200000 187.250000 ;
      RECT 0.720000 186.750000 383.200000 186.950000 ;
      RECT 0.720000 186.650000 382.480000 186.750000 ;
      RECT 0.000000 186.450000 382.480000 186.650000 ;
      RECT 0.000000 186.150000 383.200000 186.450000 ;
      RECT 0.720000 185.950000 383.200000 186.150000 ;
      RECT 0.720000 185.850000 382.480000 185.950000 ;
      RECT 0.000000 185.650000 382.480000 185.850000 ;
      RECT 0.000000 185.350000 383.200000 185.650000 ;
      RECT 0.720000 185.150000 383.200000 185.350000 ;
      RECT 0.720000 185.050000 382.480000 185.150000 ;
      RECT 0.000000 184.850000 382.480000 185.050000 ;
      RECT 0.000000 184.550000 383.200000 184.850000 ;
      RECT 0.720000 184.350000 383.200000 184.550000 ;
      RECT 0.720000 184.250000 382.480000 184.350000 ;
      RECT 0.000000 184.050000 382.480000 184.250000 ;
      RECT 0.000000 183.750000 383.200000 184.050000 ;
      RECT 0.720000 183.550000 383.200000 183.750000 ;
      RECT 0.720000 183.450000 382.480000 183.550000 ;
      RECT 0.000000 183.250000 382.480000 183.450000 ;
      RECT 0.000000 182.950000 383.200000 183.250000 ;
      RECT 0.720000 182.750000 383.200000 182.950000 ;
      RECT 0.720000 182.650000 382.480000 182.750000 ;
      RECT 0.000000 182.450000 382.480000 182.650000 ;
      RECT 0.000000 182.150000 383.200000 182.450000 ;
      RECT 0.720000 181.950000 383.200000 182.150000 ;
      RECT 0.720000 181.850000 382.480000 181.950000 ;
      RECT 0.000000 181.650000 382.480000 181.850000 ;
      RECT 0.000000 181.350000 383.200000 181.650000 ;
      RECT 0.720000 181.150000 383.200000 181.350000 ;
      RECT 0.720000 181.050000 382.480000 181.150000 ;
      RECT 0.000000 180.850000 382.480000 181.050000 ;
      RECT 0.000000 180.550000 383.200000 180.850000 ;
      RECT 0.720000 180.350000 383.200000 180.550000 ;
      RECT 0.720000 180.250000 382.480000 180.350000 ;
      RECT 0.000000 180.050000 382.480000 180.250000 ;
      RECT 0.000000 179.750000 383.200000 180.050000 ;
      RECT 0.720000 179.550000 383.200000 179.750000 ;
      RECT 0.720000 179.450000 382.480000 179.550000 ;
      RECT 0.000000 179.250000 382.480000 179.450000 ;
      RECT 0.000000 178.950000 383.200000 179.250000 ;
      RECT 0.720000 178.750000 383.200000 178.950000 ;
      RECT 0.720000 178.650000 382.480000 178.750000 ;
      RECT 0.000000 178.450000 382.480000 178.650000 ;
      RECT 0.000000 178.150000 383.200000 178.450000 ;
      RECT 0.720000 177.950000 383.200000 178.150000 ;
      RECT 0.720000 177.850000 382.480000 177.950000 ;
      RECT 0.000000 177.650000 382.480000 177.850000 ;
      RECT 0.000000 177.350000 383.200000 177.650000 ;
      RECT 0.720000 177.150000 383.200000 177.350000 ;
      RECT 0.720000 177.050000 382.480000 177.150000 ;
      RECT 0.000000 176.850000 382.480000 177.050000 ;
      RECT 0.000000 176.550000 383.200000 176.850000 ;
      RECT 0.720000 176.350000 383.200000 176.550000 ;
      RECT 0.720000 176.250000 382.480000 176.350000 ;
      RECT 0.000000 176.050000 382.480000 176.250000 ;
      RECT 0.000000 175.750000 383.200000 176.050000 ;
      RECT 0.720000 175.550000 383.200000 175.750000 ;
      RECT 0.720000 175.450000 382.480000 175.550000 ;
      RECT 0.000000 175.250000 382.480000 175.450000 ;
      RECT 0.000000 174.950000 383.200000 175.250000 ;
      RECT 0.720000 174.750000 383.200000 174.950000 ;
      RECT 0.720000 174.650000 382.480000 174.750000 ;
      RECT 0.000000 174.450000 382.480000 174.650000 ;
      RECT 0.000000 174.150000 383.200000 174.450000 ;
      RECT 0.720000 173.950000 383.200000 174.150000 ;
      RECT 0.720000 173.850000 382.480000 173.950000 ;
      RECT 0.000000 173.650000 382.480000 173.850000 ;
      RECT 0.000000 173.350000 383.200000 173.650000 ;
      RECT 0.720000 173.150000 383.200000 173.350000 ;
      RECT 0.720000 173.050000 382.480000 173.150000 ;
      RECT 0.000000 172.850000 382.480000 173.050000 ;
      RECT 0.000000 172.550000 383.200000 172.850000 ;
      RECT 0.720000 172.350000 383.200000 172.550000 ;
      RECT 0.720000 172.250000 382.480000 172.350000 ;
      RECT 0.000000 172.050000 382.480000 172.250000 ;
      RECT 0.000000 171.750000 383.200000 172.050000 ;
      RECT 0.720000 171.550000 383.200000 171.750000 ;
      RECT 0.720000 171.450000 382.480000 171.550000 ;
      RECT 0.000000 171.250000 382.480000 171.450000 ;
      RECT 0.000000 170.950000 383.200000 171.250000 ;
      RECT 0.720000 170.750000 383.200000 170.950000 ;
      RECT 0.720000 170.650000 382.480000 170.750000 ;
      RECT 0.000000 170.450000 382.480000 170.650000 ;
      RECT 0.000000 169.950000 383.200000 170.450000 ;
      RECT 0.000000 169.650000 382.480000 169.950000 ;
      RECT 0.000000 169.150000 383.200000 169.650000 ;
      RECT 0.000000 168.850000 382.480000 169.150000 ;
      RECT 0.000000 168.350000 383.200000 168.850000 ;
      RECT 0.000000 168.050000 382.480000 168.350000 ;
      RECT 0.000000 167.550000 383.200000 168.050000 ;
      RECT 0.000000 167.250000 382.480000 167.550000 ;
      RECT 0.000000 166.750000 383.200000 167.250000 ;
      RECT 0.000000 166.450000 382.480000 166.750000 ;
      RECT 0.000000 165.950000 383.200000 166.450000 ;
      RECT 0.000000 165.650000 382.480000 165.950000 ;
      RECT 0.000000 165.150000 383.200000 165.650000 ;
      RECT 0.000000 164.850000 382.480000 165.150000 ;
      RECT 0.000000 164.350000 383.200000 164.850000 ;
      RECT 0.000000 164.050000 382.480000 164.350000 ;
      RECT 0.000000 163.550000 383.200000 164.050000 ;
      RECT 0.000000 163.250000 382.480000 163.550000 ;
      RECT 0.000000 162.750000 383.200000 163.250000 ;
      RECT 0.000000 162.450000 382.480000 162.750000 ;
      RECT 0.000000 161.950000 383.200000 162.450000 ;
      RECT 0.000000 161.650000 382.480000 161.950000 ;
      RECT 0.000000 161.150000 383.200000 161.650000 ;
      RECT 0.000000 160.850000 382.480000 161.150000 ;
      RECT 0.000000 160.350000 383.200000 160.850000 ;
      RECT 0.000000 160.050000 382.480000 160.350000 ;
      RECT 0.000000 159.550000 383.200000 160.050000 ;
      RECT 0.000000 159.250000 382.480000 159.550000 ;
      RECT 0.000000 158.750000 383.200000 159.250000 ;
      RECT 0.000000 158.450000 382.480000 158.750000 ;
      RECT 0.000000 157.950000 383.200000 158.450000 ;
      RECT 0.000000 157.650000 382.480000 157.950000 ;
      RECT 0.000000 157.150000 383.200000 157.650000 ;
      RECT 0.000000 156.850000 382.480000 157.150000 ;
      RECT 0.000000 156.350000 383.200000 156.850000 ;
      RECT 0.000000 156.050000 382.480000 156.350000 ;
      RECT 0.000000 0.000000 383.200000 156.050000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 383.200000 381.800000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 383.200000 381.800000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 383.200000 381.800000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 383.200000 381.800000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 383.200000 381.800000 ;
  END
END fullchip

END LIBRARY
